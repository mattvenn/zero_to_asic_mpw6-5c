magic
tech sky130A
magscale 1 2
timestamp 1650976737
<< metal1 >>
rect 201494 703128 201500 703180
rect 201552 703168 201558 703180
rect 202782 703168 202788 703180
rect 201552 703140 202788 703168
rect 201552 703128 201558 703140
rect 202782 703128 202788 703140
rect 202840 703128 202846 703180
rect 98638 703060 98644 703112
rect 98696 703100 98702 703112
rect 332502 703100 332508 703112
rect 98696 703072 332508 703100
rect 98696 703060 98702 703072
rect 332502 703060 332508 703072
rect 332560 703060 332566 703112
rect 79318 702992 79324 703044
rect 79376 703032 79382 703044
rect 364978 703032 364984 703044
rect 79376 703004 364984 703032
rect 79376 702992 79382 703004
rect 364978 702992 364984 703004
rect 365036 702992 365042 703044
rect 106274 702924 106280 702976
rect 106332 702964 106338 702976
rect 413646 702964 413652 702976
rect 106332 702936 413652 702964
rect 106332 702924 106338 702936
rect 413646 702924 413652 702936
rect 413704 702924 413710 702976
rect 117222 702856 117228 702908
rect 117280 702896 117286 702908
rect 462314 702896 462320 702908
rect 117280 702868 462320 702896
rect 117280 702856 117286 702868
rect 462314 702856 462320 702868
rect 462372 702856 462378 702908
rect 79410 702788 79416 702840
rect 79468 702828 79474 702840
rect 429838 702828 429844 702840
rect 79468 702800 429844 702828
rect 79468 702788 79474 702800
rect 429838 702788 429844 702800
rect 429896 702788 429902 702840
rect 123478 702720 123484 702772
rect 123536 702760 123542 702772
rect 478506 702760 478512 702772
rect 123536 702732 478512 702760
rect 123536 702720 123542 702732
rect 478506 702720 478512 702732
rect 478564 702720 478570 702772
rect 119982 702652 119988 702704
rect 120040 702692 120046 702704
rect 494790 702692 494796 702704
rect 120040 702664 494796 702692
rect 120040 702652 120046 702664
rect 494790 702652 494796 702664
rect 494848 702652 494854 702704
rect 115842 702584 115848 702636
rect 115900 702624 115906 702636
rect 559650 702624 559656 702636
rect 115900 702596 559656 702624
rect 115900 702584 115906 702596
rect 559650 702584 559656 702596
rect 559708 702584 559714 702636
rect 81342 702516 81348 702568
rect 81400 702556 81406 702568
rect 527174 702556 527180 702568
rect 81400 702528 527180 702556
rect 81400 702516 81406 702528
rect 527174 702516 527180 702528
rect 527232 702516 527238 702568
rect 57238 702448 57244 702500
rect 57296 702488 57302 702500
rect 543458 702488 543464 702500
rect 57296 702460 543464 702488
rect 57296 702448 57302 702460
rect 543458 702448 543464 702460
rect 543516 702448 543522 702500
rect 86218 700340 86224 700392
rect 86276 700380 86282 700392
rect 154114 700380 154120 700392
rect 86276 700352 154120 700380
rect 86276 700340 86282 700352
rect 154114 700340 154120 700352
rect 154172 700340 154178 700392
rect 155218 700340 155224 700392
rect 155276 700380 155282 700392
rect 218974 700380 218980 700392
rect 155276 700352 218980 700380
rect 155276 700340 155282 700352
rect 218974 700340 218980 700352
rect 219032 700340 219038 700392
rect 66162 700272 66168 700324
rect 66220 700312 66226 700324
rect 170306 700312 170312 700324
rect 66220 700284 170312 700312
rect 66220 700272 66226 700284
rect 170306 700272 170312 700284
rect 170364 700272 170370 700324
rect 220078 700272 220084 700324
rect 220136 700312 220142 700324
rect 235166 700312 235172 700324
rect 220136 700284 235172 700312
rect 220136 700272 220142 700284
rect 235166 700272 235172 700284
rect 235224 700272 235230 700324
rect 341518 700272 341524 700324
rect 341576 700312 341582 700324
rect 348786 700312 348792 700324
rect 341576 700284 348792 700312
rect 341576 700272 341582 700284
rect 348786 700272 348792 700284
rect 348844 700272 348850 700324
rect 8110 700204 8116 700256
rect 8168 700244 8174 700256
rect 14458 700244 14464 700256
rect 8168 700216 14464 700244
rect 8168 700204 8174 700216
rect 14458 700204 14464 700216
rect 14516 700204 14522 700256
rect 395338 699660 395344 699712
rect 395396 699700 395402 699712
rect 397454 699700 397460 699712
rect 395396 699672 397460 699700
rect 395396 699660 395402 699672
rect 397454 699660 397460 699672
rect 397512 699660 397518 699712
rect 24302 698912 24308 698964
rect 24360 698952 24366 698964
rect 110414 698952 110420 698964
rect 24360 698924 110420 698952
rect 24360 698912 24366 698924
rect 110414 698912 110420 698924
rect 110472 698912 110478 698964
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 68278 694764 68284 694816
rect 68336 694804 68342 694816
rect 282914 694804 282920 694816
rect 68336 694776 282920 694804
rect 68336 694764 68342 694776
rect 282914 694764 282920 694776
rect 282972 694764 282978 694816
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 75178 683176 75184 683188
rect 3476 683148 75184 683176
rect 3476 683136 3482 683148
rect 75178 683136 75184 683148
rect 75236 683136 75242 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 58618 670732 58624 670744
rect 3568 670704 58624 670732
rect 3568 670692 3574 670704
rect 58618 670692 58624 670704
rect 58676 670692 58682 670744
rect 87598 670692 87604 670744
rect 87656 670732 87662 670744
rect 580166 670732 580172 670744
rect 87656 670704 580172 670732
rect 87656 670692 87662 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 35158 656928 35164 656940
rect 3476 656900 35164 656928
rect 3476 656888 3482 656900
rect 35158 656888 35164 656900
rect 35216 656888 35222 656940
rect 142798 643084 142804 643136
rect 142856 643124 142862 643136
rect 580166 643124 580172 643136
rect 142856 643096 580172 643124
rect 142856 643084 142862 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 124858 630640 124864 630692
rect 124916 630680 124922 630692
rect 579982 630680 579988 630692
rect 124916 630652 579988 630680
rect 124916 630640 124922 630652
rect 579982 630640 579988 630652
rect 580040 630640 580046 630692
rect 3510 618264 3516 618316
rect 3568 618304 3574 618316
rect 15838 618304 15844 618316
rect 3568 618276 15844 618304
rect 3568 618264 3574 618276
rect 15838 618264 15844 618276
rect 15896 618264 15902 618316
rect 3510 605820 3516 605872
rect 3568 605860 3574 605872
rect 25498 605860 25504 605872
rect 3568 605832 25504 605860
rect 3568 605820 3574 605832
rect 25498 605820 25504 605832
rect 25556 605820 25562 605872
rect 146938 590656 146944 590708
rect 146996 590696 147002 590708
rect 580166 590696 580172 590708
rect 146996 590668 580172 590696
rect 146996 590656 147002 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 32398 579680 32404 579692
rect 3384 579652 32404 579680
rect 3384 579640 3390 579652
rect 32398 579640 32404 579652
rect 32456 579640 32462 579692
rect 70302 576852 70308 576904
rect 70360 576892 70366 576904
rect 580166 576892 580172 576904
rect 70360 576864 580172 576892
rect 70360 576852 70366 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3234 565836 3240 565888
rect 3292 565876 3298 565888
rect 60734 565876 60740 565888
rect 3292 565848 60740 565876
rect 3292 565836 3298 565848
rect 60734 565836 60740 565848
rect 60792 565836 60798 565888
rect 148318 563048 148324 563100
rect 148376 563088 148382 563100
rect 580166 563088 580172 563100
rect 148376 563060 580172 563088
rect 148376 563048 148382 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 3510 553800 3516 553852
rect 3568 553840 3574 553852
rect 7558 553840 7564 553852
rect 3568 553812 7564 553840
rect 3568 553800 3574 553812
rect 7558 553800 7564 553812
rect 7616 553800 7622 553852
rect 122098 536800 122104 536852
rect 122156 536840 122162 536852
rect 579890 536840 579896 536852
rect 122156 536812 579896 536840
rect 122156 536800 122162 536812
rect 579890 536800 579896 536812
rect 579948 536800 579954 536852
rect 7558 530544 7564 530596
rect 7616 530584 7622 530596
rect 111794 530584 111800 530596
rect 7616 530556 111800 530584
rect 7616 530544 7622 530556
rect 111794 530544 111800 530556
rect 111852 530544 111858 530596
rect 2958 527144 2964 527196
rect 3016 527184 3022 527196
rect 7558 527184 7564 527196
rect 3016 527156 7564 527184
rect 3016 527144 3022 527156
rect 7558 527144 7564 527156
rect 7616 527144 7622 527196
rect 141418 524424 141424 524476
rect 141476 524464 141482 524476
rect 580166 524464 580172 524476
rect 141476 524436 580172 524464
rect 141476 524424 141482 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3510 514768 3516 514820
rect 3568 514808 3574 514820
rect 101398 514808 101404 514820
rect 3568 514780 101404 514808
rect 3568 514768 3574 514780
rect 101398 514768 101404 514780
rect 101456 514768 101462 514820
rect 76558 510620 76564 510672
rect 76616 510660 76622 510672
rect 580166 510660 580172 510672
rect 76616 510632 580172 510660
rect 76616 510620 76622 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 93118 501004 93124 501016
rect 3108 500976 93124 501004
rect 3108 500964 3114 500976
rect 93118 500964 93124 500976
rect 93176 500964 93182 501016
rect 126238 484372 126244 484424
rect 126296 484412 126302 484424
rect 580166 484412 580172 484424
rect 126296 484384 580172 484412
rect 126296 484372 126302 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 3050 474716 3056 474768
rect 3108 474756 3114 474768
rect 35250 474756 35256 474768
rect 3108 474728 35256 474756
rect 3108 474716 3114 474728
rect 35250 474716 35256 474728
rect 35308 474716 35314 474768
rect 116578 470568 116584 470620
rect 116636 470608 116642 470620
rect 580166 470608 580172 470620
rect 116636 470580 580172 470608
rect 116636 470568 116642 470580
rect 580166 470568 580172 470580
rect 580224 470568 580230 470620
rect 2774 462544 2780 462596
rect 2832 462584 2838 462596
rect 4798 462584 4804 462596
rect 2832 462556 4804 462584
rect 2832 462544 2838 462556
rect 4798 462544 4804 462556
rect 4856 462544 4862 462596
rect 97258 456764 97264 456816
rect 97316 456804 97322 456816
rect 580166 456804 580172 456816
rect 97316 456776 580172 456804
rect 97316 456764 97322 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 35158 453296 35164 453348
rect 35216 453336 35222 453348
rect 90358 453336 90364 453348
rect 35216 453308 90364 453336
rect 35216 453296 35222 453308
rect 90358 453296 90364 453308
rect 90416 453296 90422 453348
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 11698 448576 11704 448588
rect 3200 448548 11704 448576
rect 3200 448536 3206 448548
rect 11698 448536 11704 448548
rect 11756 448536 11762 448588
rect 130378 430584 130384 430636
rect 130436 430624 130442 430636
rect 579890 430624 579896 430636
rect 130436 430596 579896 430624
rect 130436 430584 130442 430596
rect 579890 430584 579896 430596
rect 579948 430584 579954 430636
rect 3510 422288 3516 422340
rect 3568 422328 3574 422340
rect 108298 422328 108304 422340
rect 3568 422300 108304 422328
rect 3568 422288 3574 422300
rect 108298 422288 108304 422300
rect 108356 422288 108362 422340
rect 72418 418140 72424 418192
rect 72476 418180 72482 418192
rect 580166 418180 580172 418192
rect 72476 418152 580172 418180
rect 72476 418140 72482 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 2866 409844 2872 409896
rect 2924 409884 2930 409896
rect 110598 409884 110604 409896
rect 2924 409856 110604 409884
rect 2924 409844 2930 409856
rect 110598 409844 110604 409856
rect 110656 409844 110662 409896
rect 97350 404336 97356 404388
rect 97408 404376 97414 404388
rect 580166 404376 580172 404388
rect 97408 404348 580172 404376
rect 97408 404336 97414 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 68830 403588 68836 403640
rect 68888 403628 68894 403640
rect 220078 403628 220084 403640
rect 68888 403600 220084 403628
rect 68888 403588 68894 403600
rect 220078 403588 220084 403600
rect 220136 403588 220142 403640
rect 15838 400868 15844 400920
rect 15896 400908 15902 400920
rect 42794 400908 42800 400920
rect 15896 400880 42800 400908
rect 15896 400868 15902 400880
rect 42794 400868 42800 400880
rect 42852 400868 42858 400920
rect 42794 400188 42800 400240
rect 42852 400228 42858 400240
rect 44082 400228 44088 400240
rect 42852 400200 44088 400228
rect 42852 400188 42858 400200
rect 44082 400188 44088 400200
rect 44140 400228 44146 400240
rect 99374 400228 99380 400240
rect 44140 400200 99380 400228
rect 44140 400188 44146 400200
rect 99374 400188 99380 400200
rect 99432 400188 99438 400240
rect 14458 399440 14464 399492
rect 14516 399480 14522 399492
rect 40862 399480 40868 399492
rect 14516 399452 40868 399480
rect 14516 399440 14522 399452
rect 40862 399440 40868 399452
rect 40920 399440 40926 399492
rect 91738 399440 91744 399492
rect 91796 399480 91802 399492
rect 97258 399480 97264 399492
rect 91796 399452 97264 399480
rect 91796 399440 91802 399452
rect 97258 399440 97264 399452
rect 97316 399440 97322 399492
rect 40862 398828 40868 398880
rect 40920 398868 40926 398880
rect 41322 398868 41328 398880
rect 40920 398840 41328 398868
rect 40920 398828 40926 398840
rect 41322 398828 41328 398840
rect 41380 398868 41386 398880
rect 89714 398868 89720 398880
rect 41380 398840 89720 398868
rect 41380 398828 41386 398840
rect 89714 398828 89720 398840
rect 89772 398828 89778 398880
rect 68738 398080 68744 398132
rect 68796 398120 68802 398132
rect 86218 398120 86224 398132
rect 68796 398092 86224 398120
rect 68796 398080 68802 398092
rect 86218 398080 86224 398092
rect 86276 398080 86282 398132
rect 3510 397468 3516 397520
rect 3568 397508 3574 397520
rect 15194 397508 15200 397520
rect 3568 397480 15200 397508
rect 3568 397468 3574 397480
rect 15194 397468 15200 397480
rect 15252 397468 15258 397520
rect 15194 396720 15200 396772
rect 15252 396760 15258 396772
rect 48222 396760 48228 396772
rect 15252 396732 48228 396760
rect 15252 396720 15258 396732
rect 48222 396720 48228 396732
rect 48280 396720 48286 396772
rect 48222 396040 48228 396092
rect 48280 396080 48286 396092
rect 111978 396080 111984 396092
rect 48280 396052 111984 396080
rect 48280 396040 48286 396052
rect 111978 396040 111984 396052
rect 112036 396040 112042 396092
rect 71038 395292 71044 395344
rect 71096 395332 71102 395344
rect 136634 395332 136640 395344
rect 71096 395304 136640 395332
rect 71096 395292 71102 395304
rect 136634 395292 136640 395304
rect 136692 395292 136698 395344
rect 135254 393932 135260 393984
rect 135312 393972 135318 393984
rect 266354 393972 266360 393984
rect 135312 393944 266360 393972
rect 135312 393932 135318 393944
rect 266354 393932 266360 393944
rect 266412 393932 266418 393984
rect 81526 393320 81532 393372
rect 81584 393360 81590 393372
rect 135254 393360 135260 393372
rect 81584 393332 135260 393360
rect 81584 393320 81590 393332
rect 135254 393320 135260 393332
rect 135312 393320 135318 393372
rect 115198 392572 115204 392624
rect 115256 392612 115262 392624
rect 299474 392612 299480 392624
rect 115256 392584 299480 392612
rect 115256 392572 115262 392584
rect 299474 392572 299480 392584
rect 299532 392572 299538 392624
rect 7558 391212 7564 391264
rect 7616 391252 7622 391264
rect 111886 391252 111892 391264
rect 7616 391224 111892 391252
rect 7616 391212 7622 391224
rect 111886 391212 111892 391224
rect 111944 391212 111950 391264
rect 118602 391212 118608 391264
rect 118660 391252 118666 391264
rect 201494 391252 201500 391264
rect 118660 391224 201500 391252
rect 118660 391212 118666 391224
rect 201494 391212 201500 391224
rect 201552 391212 201558 391264
rect 74994 390532 75000 390584
rect 75052 390572 75058 390584
rect 166258 390572 166264 390584
rect 75052 390544 166264 390572
rect 75052 390532 75058 390544
rect 166258 390532 166264 390544
rect 166316 390532 166322 390584
rect 112438 389784 112444 389836
rect 112496 389824 112502 389836
rect 148318 389824 148324 389836
rect 112496 389796 148324 389824
rect 112496 389784 112502 389796
rect 148318 389784 148324 389796
rect 148376 389784 148382 389836
rect 108298 389308 108304 389360
rect 108356 389348 108362 389360
rect 109678 389348 109684 389360
rect 108356 389320 109684 389348
rect 108356 389308 108362 389320
rect 109678 389308 109684 389320
rect 109736 389308 109742 389360
rect 65978 389240 65984 389292
rect 66036 389280 66042 389292
rect 232498 389280 232504 389292
rect 66036 389252 232504 389280
rect 66036 389240 66042 389252
rect 232498 389240 232504 389252
rect 232556 389240 232562 389292
rect 70394 389172 70400 389224
rect 70452 389212 70458 389224
rect 353294 389212 353300 389224
rect 70452 389184 353300 389212
rect 70452 389172 70458 389184
rect 353294 389172 353300 389184
rect 353352 389172 353358 389224
rect 88334 388424 88340 388476
rect 88392 388464 88398 388476
rect 117314 388464 117320 388476
rect 88392 388436 117320 388464
rect 88392 388424 88398 388436
rect 117314 388424 117320 388436
rect 117372 388424 117378 388476
rect 137094 388424 137100 388476
rect 137152 388464 137158 388476
rect 155218 388464 155224 388476
rect 137152 388436 155224 388464
rect 137152 388424 137158 388436
rect 155218 388424 155224 388436
rect 155276 388424 155282 388476
rect 102134 387880 102140 387932
rect 102192 387920 102198 387932
rect 136818 387920 136824 387932
rect 102192 387892 136824 387920
rect 102192 387880 102198 387892
rect 136818 387880 136824 387892
rect 136876 387920 136882 387932
rect 137094 387920 137100 387932
rect 136876 387892 137100 387920
rect 136876 387880 136882 387892
rect 137094 387880 137100 387892
rect 137152 387880 137158 387932
rect 85666 387812 85672 387864
rect 85724 387852 85730 387864
rect 169018 387852 169024 387864
rect 85724 387824 169024 387852
rect 85724 387812 85730 387824
rect 169018 387812 169024 387824
rect 169076 387812 169082 387864
rect 104894 387744 104900 387796
rect 104952 387784 104958 387796
rect 110690 387784 110696 387796
rect 104952 387756 110696 387784
rect 104952 387744 104958 387756
rect 110690 387744 110696 387756
rect 110748 387744 110754 387796
rect 40034 387064 40040 387116
rect 40092 387104 40098 387116
rect 51074 387104 51080 387116
rect 40092 387076 51080 387104
rect 40092 387064 40098 387076
rect 51074 387064 51080 387076
rect 51132 387064 51138 387116
rect 76650 387064 76656 387116
rect 76708 387104 76714 387116
rect 97350 387104 97356 387116
rect 76708 387076 97356 387104
rect 76708 387064 76714 387076
rect 97350 387064 97356 387076
rect 97408 387064 97414 387116
rect 113910 387064 113916 387116
rect 113968 387104 113974 387116
rect 580258 387104 580264 387116
rect 113968 387076 580264 387104
rect 113968 387064 113974 387076
rect 580258 387064 580264 387076
rect 580316 387064 580322 387116
rect 51074 386520 51080 386572
rect 51132 386560 51138 386572
rect 52362 386560 52368 386572
rect 51132 386532 52368 386560
rect 51132 386520 51138 386532
rect 52362 386520 52368 386532
rect 52420 386560 52426 386572
rect 76742 386560 76748 386572
rect 52420 386532 76748 386560
rect 52420 386520 52426 386532
rect 76742 386520 76748 386532
rect 76800 386520 76806 386572
rect 100754 386520 100760 386572
rect 100812 386560 100818 386572
rect 101398 386560 101404 386572
rect 100812 386532 101404 386560
rect 100812 386520 100818 386532
rect 101398 386520 101404 386532
rect 101456 386560 101462 386572
rect 147674 386560 147680 386572
rect 101456 386532 147680 386560
rect 101456 386520 101462 386532
rect 147674 386520 147680 386532
rect 147732 386520 147738 386572
rect 68830 386452 68836 386504
rect 68888 386492 68894 386504
rect 132494 386492 132500 386504
rect 68888 386464 132500 386492
rect 68888 386452 68894 386464
rect 132494 386452 132500 386464
rect 132552 386452 132558 386504
rect 73706 386384 73712 386436
rect 73764 386424 73770 386436
rect 313918 386424 313924 386436
rect 73764 386396 313924 386424
rect 73764 386384 73770 386396
rect 313918 386384 313924 386396
rect 313976 386384 313982 386436
rect 84930 386316 84936 386368
rect 84988 386356 84994 386368
rect 87598 386356 87604 386368
rect 84988 386328 87604 386356
rect 84988 386316 84994 386328
rect 87598 386316 87604 386328
rect 87656 386316 87662 386368
rect 109678 385364 109684 385416
rect 109736 385404 109742 385416
rect 124214 385404 124220 385416
rect 109736 385376 124220 385404
rect 109736 385364 109742 385376
rect 124214 385364 124220 385376
rect 124272 385364 124278 385416
rect 88242 385296 88248 385348
rect 88300 385336 88306 385348
rect 121454 385336 121460 385348
rect 88300 385308 121460 385336
rect 88300 385296 88306 385308
rect 121454 385296 121460 385308
rect 121512 385296 121518 385348
rect 90358 385228 90364 385280
rect 90416 385268 90422 385280
rect 125594 385268 125600 385280
rect 90416 385240 125600 385268
rect 90416 385228 90422 385240
rect 125594 385228 125600 385240
rect 125652 385228 125658 385280
rect 81342 385160 81348 385212
rect 81400 385200 81406 385212
rect 128538 385200 128544 385212
rect 81400 385172 128544 385200
rect 81400 385160 81406 385172
rect 128538 385160 128544 385172
rect 128596 385160 128602 385212
rect 57790 385092 57796 385144
rect 57848 385132 57854 385144
rect 98638 385132 98644 385144
rect 57848 385104 98644 385132
rect 57848 385092 57854 385104
rect 98638 385092 98644 385104
rect 98696 385092 98702 385144
rect 100662 385092 100668 385144
rect 100720 385132 100726 385144
rect 160738 385132 160744 385144
rect 100720 385104 160744 385132
rect 100720 385092 100726 385104
rect 160738 385092 160744 385104
rect 160796 385092 160802 385144
rect 70210 385024 70216 385076
rect 70268 385064 70274 385076
rect 76558 385064 76564 385076
rect 70268 385036 76564 385064
rect 70268 385024 70274 385036
rect 76558 385024 76564 385036
rect 76616 385024 76622 385076
rect 94590 385024 94596 385076
rect 94648 385064 94654 385076
rect 309778 385064 309784 385076
rect 94648 385036 309784 385064
rect 94648 385024 94654 385036
rect 309778 385024 309784 385036
rect 309836 385024 309842 385076
rect 68370 384140 68376 384192
rect 68428 384180 68434 384192
rect 72418 384180 72424 384192
rect 68428 384152 72424 384180
rect 68428 384140 68434 384152
rect 72418 384140 72424 384152
rect 72476 384140 72482 384192
rect 96522 383936 96528 383988
rect 96580 383976 96586 383988
rect 128354 383976 128360 383988
rect 96580 383948 128360 383976
rect 96580 383936 96586 383948
rect 128354 383936 128360 383948
rect 128412 383936 128418 383988
rect 93118 383868 93124 383920
rect 93176 383908 93182 383920
rect 132586 383908 132592 383920
rect 93176 383880 132592 383908
rect 93176 383868 93182 383880
rect 132586 383868 132592 383880
rect 132644 383868 132650 383920
rect 73062 383800 73068 383852
rect 73120 383840 73126 383852
rect 118694 383840 118700 383852
rect 73120 383812 118700 383840
rect 73120 383800 73126 383812
rect 118694 383800 118700 383812
rect 118752 383800 118758 383852
rect 49602 383732 49608 383784
rect 49660 383772 49666 383784
rect 71038 383772 71044 383784
rect 49660 383744 71044 383772
rect 49660 383732 49666 383744
rect 71038 383732 71044 383744
rect 71096 383732 71102 383784
rect 97902 383732 97908 383784
rect 97960 383772 97966 383784
rect 195238 383772 195244 383784
rect 97960 383744 195244 383772
rect 97960 383732 97966 383744
rect 195238 383732 195244 383744
rect 195296 383732 195302 383784
rect 62022 383664 62028 383716
rect 62080 383704 62086 383716
rect 84930 383704 84936 383716
rect 62080 383676 84936 383704
rect 62080 383664 62086 383676
rect 84930 383664 84936 383676
rect 84988 383664 84994 383716
rect 103882 383664 103888 383716
rect 103940 383704 103946 383716
rect 215938 383704 215944 383716
rect 103940 383676 215944 383704
rect 103940 383664 103946 383676
rect 215938 383664 215944 383676
rect 215996 383664 216002 383716
rect 84562 382916 84568 382968
rect 84620 382956 84626 382968
rect 100662 382956 100668 382968
rect 84620 382928 100668 382956
rect 84620 382916 84626 382928
rect 100662 382916 100668 382928
rect 100720 382916 100726 382968
rect 101858 382644 101864 382696
rect 101916 382684 101922 382696
rect 209038 382684 209044 382696
rect 101916 382656 209044 382684
rect 101916 382644 101922 382656
rect 209038 382644 209044 382656
rect 209096 382644 209102 382696
rect 77846 382576 77852 382628
rect 77904 382616 77910 382628
rect 79410 382616 79416 382628
rect 77904 382588 79416 382616
rect 77904 382576 77910 382588
rect 79410 382576 79416 382588
rect 79468 382576 79474 382628
rect 96154 382576 96160 382628
rect 96212 382616 96218 382628
rect 280798 382616 280804 382628
rect 96212 382588 280804 382616
rect 96212 382576 96218 382588
rect 280798 382576 280804 382588
rect 280856 382576 280862 382628
rect 59262 382508 59268 382560
rect 59320 382548 59326 382560
rect 70210 382548 70216 382560
rect 59320 382520 70216 382548
rect 59320 382508 59326 382520
rect 70210 382508 70216 382520
rect 70268 382508 70274 382560
rect 76650 382548 76656 382560
rect 70366 382520 76656 382548
rect 60642 382440 60648 382492
rect 60700 382480 60706 382492
rect 70366 382480 70394 382520
rect 76650 382508 76656 382520
rect 76708 382508 76714 382560
rect 87690 382508 87696 382560
rect 87748 382548 87754 382560
rect 109862 382548 109868 382560
rect 87748 382520 109868 382548
rect 87748 382508 87754 382520
rect 109862 382508 109868 382520
rect 109920 382508 109926 382560
rect 77846 382480 77852 382492
rect 60700 382452 70394 382480
rect 74736 382452 77852 382480
rect 60700 382440 60706 382452
rect 55122 382372 55128 382424
rect 55180 382412 55186 382424
rect 74736 382412 74764 382452
rect 77846 382440 77852 382452
rect 77904 382440 77910 382492
rect 80698 382440 80704 382492
rect 80756 382480 80762 382492
rect 106826 382480 106832 382492
rect 80756 382452 106832 382480
rect 80756 382440 80762 382452
rect 106826 382440 106832 382452
rect 106884 382440 106890 382492
rect 55180 382384 74764 382412
rect 55180 382372 55186 382384
rect 74810 382372 74816 382424
rect 74868 382412 74874 382424
rect 89806 382412 89812 382424
rect 74868 382384 89812 382412
rect 74868 382372 74874 382384
rect 89806 382372 89812 382384
rect 89864 382372 89870 382424
rect 92842 382372 92848 382424
rect 92900 382412 92906 382424
rect 133966 382412 133972 382424
rect 92900 382384 133972 382412
rect 92900 382372 92906 382384
rect 133966 382372 133972 382384
rect 134024 382372 134030 382424
rect 56410 382304 56416 382356
rect 56468 382344 56474 382356
rect 81894 382344 81900 382356
rect 56468 382316 81900 382344
rect 56468 382304 56474 382316
rect 81894 382304 81900 382316
rect 81952 382304 81958 382356
rect 85298 382304 85304 382356
rect 85356 382344 85362 382356
rect 104802 382344 104808 382356
rect 85356 382316 104808 382344
rect 85356 382304 85362 382316
rect 104802 382304 104808 382316
rect 104860 382304 104866 382356
rect 21358 382236 21364 382288
rect 21416 382276 21422 382288
rect 72050 382276 72056 382288
rect 21416 382248 72056 382276
rect 21416 382236 21422 382248
rect 72050 382236 72056 382248
rect 72108 382276 72114 382288
rect 73062 382276 73068 382288
rect 72108 382248 73068 382276
rect 72108 382236 72114 382248
rect 73062 382236 73068 382248
rect 73120 382236 73126 382288
rect 106182 382236 106188 382288
rect 106240 382276 106246 382288
rect 113818 382276 113824 382288
rect 106240 382248 113824 382276
rect 106240 382236 106246 382248
rect 113818 382236 113824 382248
rect 113876 382236 113882 382288
rect 74902 382168 74908 382220
rect 74960 382208 74966 382220
rect 75178 382208 75184 382220
rect 74960 382180 75184 382208
rect 74960 382168 74966 382180
rect 75178 382168 75184 382180
rect 75236 382168 75242 382220
rect 97442 381080 97448 381132
rect 97500 381120 97506 381132
rect 109770 381120 109776 381132
rect 97500 381092 109776 381120
rect 97500 381080 97506 381092
rect 109770 381080 109776 381092
rect 109828 381080 109834 381132
rect 50982 381012 50988 381064
rect 51040 381052 51046 381064
rect 79318 381052 79324 381064
rect 51040 381024 79324 381052
rect 51040 381012 51046 381024
rect 79318 381012 79324 381024
rect 79376 381012 79382 381064
rect 104618 381012 104624 381064
rect 104676 381052 104682 381064
rect 136634 381052 136640 381064
rect 104676 381024 136640 381052
rect 104676 381012 104682 381024
rect 136634 381012 136640 381024
rect 136692 381012 136698 381064
rect 74902 380944 74908 380996
rect 74960 380984 74966 380996
rect 122834 380984 122840 380996
rect 74960 380956 122840 380984
rect 74960 380944 74966 380956
rect 122834 380944 122840 380956
rect 122892 380944 122898 380996
rect 50890 380876 50896 380928
rect 50948 380916 50954 380928
rect 111794 380916 111800 380928
rect 50948 380888 111800 380916
rect 50948 380876 50954 380888
rect 111794 380876 111800 380888
rect 111852 380916 111858 380928
rect 112162 380916 112168 380928
rect 111852 380888 112168 380916
rect 111852 380876 111858 380888
rect 112162 380876 112168 380888
rect 112220 380876 112226 380928
rect 106826 380196 106832 380248
rect 106884 380236 106890 380248
rect 131206 380236 131212 380248
rect 106884 380208 131212 380236
rect 106884 380196 106890 380208
rect 131206 380196 131212 380208
rect 131264 380196 131270 380248
rect 104802 380128 104808 380180
rect 104860 380168 104866 380180
rect 173158 380168 173164 380180
rect 104860 380140 173164 380168
rect 104860 380128 104866 380140
rect 173158 380128 173164 380140
rect 173216 380128 173222 380180
rect 66070 380060 66076 380112
rect 66128 380100 66134 380112
rect 71958 380100 71964 380112
rect 66128 380072 71964 380100
rect 66128 380060 66134 380072
rect 71958 380060 71964 380072
rect 72016 380060 72022 380112
rect 71682 379720 71688 379772
rect 71740 379760 71746 379772
rect 109494 379760 109500 379772
rect 71740 379732 109500 379760
rect 71740 379720 71746 379732
rect 109494 379720 109500 379732
rect 109552 379720 109558 379772
rect 34330 379652 34336 379704
rect 34388 379692 34394 379704
rect 78766 379692 78772 379704
rect 34388 379664 78772 379692
rect 34388 379652 34394 379664
rect 78766 379652 78772 379664
rect 78824 379652 78830 379704
rect 53650 379584 53656 379636
rect 53708 379624 53714 379636
rect 99926 379624 99932 379636
rect 53708 379596 99932 379624
rect 53708 379584 53714 379596
rect 99926 379584 99932 379596
rect 99984 379584 99990 379636
rect 103146 379584 103152 379636
rect 103204 379624 103210 379636
rect 121546 379624 121552 379636
rect 103204 379596 121552 379624
rect 103204 379584 103210 379596
rect 121546 379584 121552 379596
rect 121604 379584 121610 379636
rect 43990 379516 43996 379568
rect 44048 379556 44054 379568
rect 105078 379556 105084 379568
rect 44048 379528 105084 379556
rect 44048 379516 44054 379528
rect 105078 379516 105084 379528
rect 105136 379516 105142 379568
rect 107010 379516 107016 379568
rect 107068 379556 107074 379568
rect 114646 379556 114652 379568
rect 107068 379528 114652 379556
rect 107068 379516 107074 379528
rect 114646 379516 114652 379528
rect 114704 379516 114710 379568
rect 107654 379448 107660 379500
rect 107712 379488 107718 379500
rect 109678 379488 109684 379500
rect 107712 379460 109684 379488
rect 107712 379448 107718 379460
rect 109678 379448 109684 379460
rect 109736 379448 109742 379500
rect 71682 379380 71688 379432
rect 71740 379420 71746 379432
rect 73706 379420 73712 379432
rect 71740 379392 73712 379420
rect 71740 379380 71746 379392
rect 73706 379380 73712 379392
rect 73764 379380 73770 379432
rect 108298 379244 108304 379296
rect 108356 379284 108362 379296
rect 108356 379256 122834 379284
rect 108356 379244 108362 379256
rect 111794 378428 111800 378480
rect 111852 378468 111858 378480
rect 114002 378468 114008 378480
rect 111852 378440 114008 378468
rect 111852 378428 111858 378440
rect 114002 378428 114008 378440
rect 114060 378428 114066 378480
rect 122806 378196 122834 379256
rect 140774 378196 140780 378208
rect 122806 378168 140780 378196
rect 140774 378156 140780 378168
rect 140832 378156 140838 378208
rect 39942 376796 39948 376848
rect 40000 376836 40006 376848
rect 67634 376836 67640 376848
rect 40000 376808 67640 376836
rect 40000 376796 40006 376808
rect 67634 376796 67640 376808
rect 67692 376796 67698 376848
rect 111794 376796 111800 376848
rect 111852 376836 111858 376848
rect 119338 376836 119344 376848
rect 111852 376808 119344 376836
rect 111852 376796 111858 376808
rect 119338 376796 119344 376808
rect 119396 376796 119402 376848
rect 35802 376728 35808 376780
rect 35860 376768 35866 376780
rect 67726 376768 67732 376780
rect 35860 376740 67732 376768
rect 35860 376728 35866 376740
rect 67726 376728 67732 376740
rect 67784 376728 67790 376780
rect 115750 376728 115756 376780
rect 115808 376768 115814 376780
rect 128446 376768 128452 376780
rect 115808 376740 128452 376768
rect 115808 376728 115814 376740
rect 128446 376728 128452 376740
rect 128504 376728 128510 376780
rect 111794 375708 111800 375760
rect 111852 375748 111858 375760
rect 115750 375748 115756 375760
rect 111852 375720 115756 375748
rect 111852 375708 111858 375720
rect 115750 375708 115756 375720
rect 115808 375708 115814 375760
rect 64782 375368 64788 375420
rect 64840 375408 64846 375420
rect 67634 375408 67640 375420
rect 64840 375380 67640 375408
rect 64840 375368 64846 375380
rect 67634 375368 67640 375380
rect 67692 375368 67698 375420
rect 112070 375368 112076 375420
rect 112128 375408 112134 375420
rect 116670 375408 116676 375420
rect 112128 375380 116676 375408
rect 112128 375368 112134 375380
rect 116670 375368 116676 375380
rect 116728 375368 116734 375420
rect 3510 374620 3516 374672
rect 3568 374660 3574 374672
rect 67542 374660 67548 374672
rect 3568 374632 67548 374660
rect 3568 374620 3574 374632
rect 67542 374620 67548 374632
rect 67600 374620 67606 374672
rect 53742 374008 53748 374060
rect 53800 374048 53806 374060
rect 57238 374048 57244 374060
rect 53800 374020 57244 374048
rect 53800 374008 53806 374020
rect 57238 374008 57244 374020
rect 57296 374048 57302 374060
rect 57296 374020 57974 374048
rect 57296 374008 57302 374020
rect 57946 373980 57974 374020
rect 111794 374008 111800 374060
rect 111852 374048 111858 374060
rect 196618 374048 196624 374060
rect 111852 374020 196624 374048
rect 111852 374008 111858 374020
rect 196618 374008 196624 374020
rect 196676 374008 196682 374060
rect 67634 373980 67640 373992
rect 57946 373952 67640 373980
rect 67634 373940 67640 373952
rect 67692 373940 67698 373992
rect 114002 373260 114008 373312
rect 114060 373300 114066 373312
rect 349154 373300 349160 373312
rect 114060 373272 349160 373300
rect 114060 373260 114066 373272
rect 349154 373260 349160 373272
rect 349212 373260 349218 373312
rect 111978 372784 111984 372836
rect 112036 372824 112042 372836
rect 112162 372824 112168 372836
rect 112036 372796 112168 372824
rect 112036 372784 112042 372796
rect 112162 372784 112168 372796
rect 112220 372784 112226 372836
rect 65978 372512 65984 372564
rect 66036 372552 66042 372564
rect 67634 372552 67640 372564
rect 66036 372524 67640 372552
rect 66036 372512 66042 372524
rect 67634 372512 67640 372524
rect 67692 372512 67698 372564
rect 112346 372512 112352 372564
rect 112404 372552 112410 372564
rect 113910 372552 113916 372564
rect 112404 372524 113916 372552
rect 112404 372512 112410 372524
rect 113910 372512 113916 372524
rect 113968 372512 113974 372564
rect 3326 371220 3332 371272
rect 3384 371260 3390 371272
rect 39298 371260 39304 371272
rect 3384 371232 39304 371260
rect 3384 371220 3390 371232
rect 39298 371220 39304 371232
rect 39356 371220 39362 371272
rect 67266 371220 67272 371272
rect 67324 371260 67330 371272
rect 68646 371260 68652 371272
rect 67324 371232 68652 371260
rect 67324 371220 67330 371232
rect 68646 371220 68652 371232
rect 68704 371220 68710 371272
rect 109678 370472 109684 370524
rect 109736 370512 109742 370524
rect 271874 370512 271880 370524
rect 109736 370484 271880 370512
rect 109736 370472 109742 370484
rect 271874 370472 271880 370484
rect 271932 370472 271938 370524
rect 111794 369928 111800 369980
rect 111852 369968 111858 369980
rect 114462 369968 114468 369980
rect 111852 369940 114468 369968
rect 111852 369928 111858 369940
rect 114462 369928 114468 369940
rect 114520 369928 114526 369980
rect 112346 369112 112352 369164
rect 112404 369152 112410 369164
rect 120074 369152 120080 369164
rect 112404 369124 120080 369152
rect 112404 369112 112410 369124
rect 120074 369112 120080 369124
rect 120132 369112 120138 369164
rect 60458 368500 60464 368552
rect 60516 368540 60522 368552
rect 67634 368540 67640 368552
rect 60516 368512 67640 368540
rect 60516 368500 60522 368512
rect 67634 368500 67640 368512
rect 67692 368500 67698 368552
rect 37182 367072 37188 367124
rect 37240 367112 37246 367124
rect 67634 367112 67640 367124
rect 37240 367084 67640 367112
rect 37240 367072 37246 367084
rect 67634 367072 67640 367084
rect 67692 367072 67698 367124
rect 111794 367072 111800 367124
rect 111852 367112 111858 367124
rect 324958 367112 324964 367124
rect 111852 367084 324964 367112
rect 111852 367072 111858 367084
rect 324958 367072 324964 367084
rect 325016 367072 325022 367124
rect 63402 365712 63408 365764
rect 63460 365752 63466 365764
rect 67634 365752 67640 365764
rect 63460 365724 67640 365752
rect 63460 365712 63466 365724
rect 67634 365712 67640 365724
rect 67692 365712 67698 365764
rect 109310 365712 109316 365764
rect 109368 365752 109374 365764
rect 110322 365752 110328 365764
rect 109368 365724 110328 365752
rect 109368 365712 109374 365724
rect 110322 365712 110328 365724
rect 110380 365752 110386 365764
rect 118602 365752 118608 365764
rect 110380 365724 118608 365752
rect 110380 365712 110386 365724
rect 118602 365712 118608 365724
rect 118660 365712 118666 365764
rect 111794 364760 111800 364812
rect 111852 364800 111858 364812
rect 114554 364800 114560 364812
rect 111852 364772 114560 364800
rect 111852 364760 111858 364772
rect 114554 364760 114560 364772
rect 114612 364760 114618 364812
rect 111794 364624 111800 364676
rect 111852 364664 111858 364676
rect 112070 364664 112076 364676
rect 111852 364636 112076 364664
rect 111852 364624 111858 364636
rect 112070 364624 112076 364636
rect 112128 364624 112134 364676
rect 63310 364420 63316 364472
rect 63368 364460 63374 364472
rect 67634 364460 67640 364472
rect 63368 364432 67640 364460
rect 63368 364420 63374 364432
rect 67634 364420 67640 364432
rect 67692 364420 67698 364472
rect 59170 364352 59176 364404
rect 59228 364392 59234 364404
rect 67726 364392 67732 364404
rect 59228 364364 67732 364392
rect 59228 364352 59234 364364
rect 67726 364352 67732 364364
rect 67784 364352 67790 364404
rect 111978 364352 111984 364404
rect 112036 364392 112042 364404
rect 142154 364392 142160 364404
rect 112036 364364 142160 364392
rect 112036 364352 112042 364364
rect 142154 364352 142160 364364
rect 142212 364352 142218 364404
rect 316770 364352 316776 364404
rect 316828 364392 316834 364404
rect 579614 364392 579620 364404
rect 316828 364364 579620 364392
rect 316828 364352 316834 364364
rect 579614 364352 579620 364364
rect 579672 364352 579678 364404
rect 119338 363604 119344 363656
rect 119396 363644 119402 363656
rect 282914 363644 282920 363656
rect 119396 363616 282920 363644
rect 119396 363604 119402 363616
rect 282914 363604 282920 363616
rect 282972 363604 282978 363656
rect 111886 362244 111892 362296
rect 111944 362284 111950 362296
rect 122098 362284 122104 362296
rect 111944 362256 122104 362284
rect 111944 362244 111950 362256
rect 122098 362244 122104 362256
rect 122156 362244 122162 362296
rect 111978 362176 111984 362228
rect 112036 362216 112042 362228
rect 116578 362216 116584 362228
rect 112036 362188 116584 362216
rect 112036 362176 112042 362188
rect 116578 362176 116584 362188
rect 116636 362176 116642 362228
rect 118602 362176 118608 362228
rect 118660 362216 118666 362228
rect 580350 362216 580356 362228
rect 118660 362188 580356 362216
rect 118660 362176 118666 362188
rect 580350 362176 580356 362188
rect 580408 362176 580414 362228
rect 34422 361564 34428 361616
rect 34480 361604 34486 361616
rect 67634 361604 67640 361616
rect 34480 361576 67640 361604
rect 34480 361564 34486 361576
rect 67634 361564 67640 361576
rect 67692 361564 67698 361616
rect 109586 361496 109592 361548
rect 109644 361536 109650 361548
rect 123478 361536 123484 361548
rect 109644 361508 123484 361536
rect 109644 361496 109650 361508
rect 123478 361496 123484 361508
rect 123536 361496 123542 361548
rect 61838 360272 61844 360324
rect 61896 360312 61902 360324
rect 67726 360312 67732 360324
rect 61896 360284 67732 360312
rect 61896 360272 61902 360284
rect 67726 360272 67732 360284
rect 67784 360312 67790 360324
rect 68278 360312 68284 360324
rect 67784 360284 68284 360312
rect 67784 360272 67790 360284
rect 68278 360272 68284 360284
rect 68336 360272 68342 360324
rect 111886 360272 111892 360324
rect 111944 360312 111950 360324
rect 202138 360312 202144 360324
rect 111944 360284 202144 360312
rect 111944 360272 111950 360284
rect 202138 360272 202144 360284
rect 202196 360272 202202 360324
rect 48130 360204 48136 360256
rect 48188 360244 48194 360256
rect 67634 360244 67640 360256
rect 48188 360216 67640 360244
rect 48188 360204 48194 360216
rect 67634 360204 67640 360216
rect 67692 360204 67698 360256
rect 111886 358844 111892 358896
rect 111944 358884 111950 358896
rect 122926 358884 122932 358896
rect 111944 358856 122932 358884
rect 111944 358844 111950 358856
rect 122926 358844 122932 358856
rect 122984 358844 122990 358896
rect 37090 358776 37096 358828
rect 37148 358816 37154 358828
rect 67634 358816 67640 358828
rect 37148 358788 67640 358816
rect 37148 358776 37154 358788
rect 67634 358776 67640 358788
rect 67692 358776 67698 358828
rect 111978 358776 111984 358828
rect 112036 358816 112042 358828
rect 186958 358816 186964 358828
rect 112036 358788 186964 358816
rect 112036 358776 112042 358788
rect 186958 358776 186964 358788
rect 187016 358776 187022 358828
rect 57882 357484 57888 357536
rect 57940 357524 57946 357536
rect 67726 357524 67732 357536
rect 57940 357496 67732 357524
rect 57940 357484 57946 357496
rect 67726 357484 67732 357496
rect 67784 357484 67790 357536
rect 3326 357416 3332 357468
rect 3384 357456 3390 357468
rect 22738 357456 22744 357468
rect 3384 357428 22744 357456
rect 3384 357416 3390 357428
rect 22738 357416 22744 357428
rect 22796 357416 22802 357468
rect 56502 357416 56508 357468
rect 56560 357456 56566 357468
rect 67634 357456 67640 357468
rect 56560 357428 67640 357456
rect 56560 357416 56566 357428
rect 67634 357416 67640 357428
rect 67692 357416 67698 357468
rect 118510 357456 118516 357468
rect 118160 357428 118516 357456
rect 111886 357348 111892 357400
rect 111944 357388 111950 357400
rect 118160 357388 118188 357428
rect 118510 357416 118516 357428
rect 118568 357456 118574 357468
rect 127066 357456 127072 357468
rect 118568 357428 127072 357456
rect 118568 357416 118574 357428
rect 127066 357416 127072 357428
rect 127124 357416 127130 357468
rect 111944 357360 118188 357388
rect 111944 357348 111950 357360
rect 55030 356056 55036 356108
rect 55088 356096 55094 356108
rect 67634 356096 67640 356108
rect 55088 356068 67640 356096
rect 55088 356056 55094 356068
rect 67634 356056 67640 356068
rect 67692 356056 67698 356108
rect 111886 356056 111892 356108
rect 111944 356096 111950 356108
rect 211798 356096 211804 356108
rect 111944 356068 211804 356096
rect 111944 356056 111950 356068
rect 211798 356056 211804 356068
rect 211856 356056 211862 356108
rect 60550 354764 60556 354816
rect 60608 354804 60614 354816
rect 66162 354804 66168 354816
rect 60608 354776 66168 354804
rect 60608 354764 60614 354776
rect 66162 354764 66168 354776
rect 66220 354804 66226 354816
rect 67726 354804 67732 354816
rect 66220 354776 67732 354804
rect 66220 354764 66226 354776
rect 67726 354764 67732 354776
rect 67784 354764 67790 354816
rect 64598 354696 64604 354748
rect 64656 354736 64662 354748
rect 67634 354736 67640 354748
rect 64656 354708 67640 354736
rect 64656 354696 64662 354708
rect 67634 354696 67640 354708
rect 67692 354696 67698 354748
rect 111886 354696 111892 354748
rect 111944 354736 111950 354748
rect 206278 354736 206284 354748
rect 111944 354708 206284 354736
rect 111944 354696 111950 354708
rect 206278 354696 206284 354708
rect 206336 354696 206342 354748
rect 65978 353336 65984 353388
rect 66036 353376 66042 353388
rect 68094 353376 68100 353388
rect 66036 353348 68100 353376
rect 66036 353336 66042 353348
rect 68094 353336 68100 353348
rect 68152 353336 68158 353388
rect 46842 353268 46848 353320
rect 46900 353308 46906 353320
rect 67634 353308 67640 353320
rect 46900 353280 67640 353308
rect 46900 353268 46906 353280
rect 67634 353268 67640 353280
rect 67692 353268 67698 353320
rect 111886 353268 111892 353320
rect 111944 353308 111950 353320
rect 139394 353308 139400 353320
rect 111944 353280 139400 353308
rect 111944 353268 111950 353280
rect 139394 353268 139400 353280
rect 139452 353268 139458 353320
rect 61930 351908 61936 351960
rect 61988 351948 61994 351960
rect 67634 351948 67640 351960
rect 61988 351920 67640 351948
rect 61988 351908 61994 351920
rect 67634 351908 67640 351920
rect 67692 351908 67698 351960
rect 111058 351908 111064 351960
rect 111116 351948 111122 351960
rect 129734 351948 129740 351960
rect 111116 351920 129740 351948
rect 111116 351908 111122 351920
rect 129734 351908 129740 351920
rect 129792 351908 129798 351960
rect 42702 350548 42708 350600
rect 42760 350588 42766 350600
rect 67634 350588 67640 350600
rect 42760 350560 67640 350588
rect 42760 350548 42766 350560
rect 67634 350548 67640 350560
rect 67692 350548 67698 350600
rect 111886 350548 111892 350600
rect 111944 350588 111950 350600
rect 143534 350588 143540 350600
rect 111944 350560 143540 350588
rect 111944 350548 111950 350560
rect 143534 350548 143540 350560
rect 143592 350588 143598 350600
rect 146938 350588 146944 350600
rect 143592 350560 146944 350588
rect 143592 350548 143598 350560
rect 146938 350548 146944 350560
rect 146996 350548 147002 350600
rect 112162 349188 112168 349240
rect 112220 349228 112226 349240
rect 135162 349228 135168 349240
rect 112220 349200 135168 349228
rect 112220 349188 112226 349200
rect 135162 349188 135168 349200
rect 135220 349188 135226 349240
rect 111886 349120 111892 349172
rect 111944 349160 111950 349172
rect 269758 349160 269764 349172
rect 111944 349132 269764 349160
rect 111944 349120 111950 349132
rect 269758 349120 269764 349132
rect 269816 349120 269822 349172
rect 135162 348372 135168 348424
rect 135220 348412 135226 348424
rect 346394 348412 346400 348424
rect 135220 348384 346400 348412
rect 135220 348372 135226 348384
rect 346394 348372 346400 348384
rect 346452 348372 346458 348424
rect 64690 347828 64696 347880
rect 64748 347868 64754 347880
rect 67634 347868 67640 347880
rect 64748 347840 67640 347868
rect 64748 347828 64754 347840
rect 67634 347828 67640 347840
rect 67692 347828 67698 347880
rect 45462 347760 45468 347812
rect 45520 347800 45526 347812
rect 67726 347800 67732 347812
rect 45520 347772 67732 347800
rect 45520 347760 45526 347772
rect 67726 347760 67732 347772
rect 67784 347760 67790 347812
rect 111886 347760 111892 347812
rect 111944 347800 111950 347812
rect 206370 347800 206376 347812
rect 111944 347772 206376 347800
rect 111944 347760 111950 347772
rect 206370 347760 206376 347772
rect 206428 347760 206434 347812
rect 111886 346400 111892 346452
rect 111944 346440 111950 346452
rect 278038 346440 278044 346452
rect 111944 346412 278044 346440
rect 111944 346400 111950 346412
rect 278038 346400 278044 346412
rect 278096 346400 278102 346452
rect 3326 346332 3332 346384
rect 3384 346372 3390 346384
rect 21358 346372 21364 346384
rect 3384 346344 21364 346372
rect 3384 346332 3390 346344
rect 21358 346332 21364 346344
rect 21416 346332 21422 346384
rect 111886 345108 111892 345160
rect 111944 345148 111950 345160
rect 123018 345148 123024 345160
rect 111944 345120 123024 345148
rect 111944 345108 111950 345120
rect 123018 345108 123024 345120
rect 123076 345108 123082 345160
rect 112162 345040 112168 345092
rect 112220 345080 112226 345092
rect 216030 345080 216036 345092
rect 112220 345052 216036 345080
rect 112220 345040 112226 345052
rect 216030 345040 216036 345052
rect 216088 345040 216094 345092
rect 60734 344972 60740 345024
rect 60792 345012 60798 345024
rect 67634 345012 67640 345024
rect 60792 344984 67640 345012
rect 60792 344972 60798 344984
rect 67634 344972 67640 344984
rect 67692 344972 67698 345024
rect 22738 344292 22744 344344
rect 22796 344332 22802 344344
rect 51074 344332 51080 344344
rect 22796 344304 51080 344332
rect 22796 344292 22802 344304
rect 51074 344292 51080 344304
rect 51132 344292 51138 344344
rect 54938 344292 54944 344344
rect 54996 344332 55002 344344
rect 60734 344332 60740 344344
rect 54996 344304 60740 344332
rect 54996 344292 55002 344304
rect 60734 344292 60740 344304
rect 60792 344292 60798 344344
rect 111978 344224 111984 344276
rect 112036 344264 112042 344276
rect 112162 344264 112168 344276
rect 112036 344236 112168 344264
rect 112036 344224 112042 344236
rect 112162 344224 112168 344236
rect 112220 344224 112226 344276
rect 111886 343816 111892 343868
rect 111944 343856 111950 343868
rect 115842 343856 115848 343868
rect 111944 343828 115848 343856
rect 111944 343816 111950 343828
rect 115842 343816 115848 343828
rect 115900 343816 115906 343868
rect 51074 343612 51080 343664
rect 51132 343652 51138 343664
rect 52178 343652 52184 343664
rect 51132 343624 52184 343652
rect 51132 343612 51138 343624
rect 52178 343612 52184 343624
rect 52236 343652 52242 343664
rect 67726 343652 67732 343664
rect 52236 343624 67732 343652
rect 52236 343612 52242 343624
rect 67726 343612 67732 343624
rect 67784 343612 67790 343664
rect 111978 343612 111984 343664
rect 112036 343652 112042 343664
rect 316678 343652 316684 343664
rect 112036 343624 316684 343652
rect 112036 343612 112042 343624
rect 316678 343612 316684 343624
rect 316736 343612 316742 343664
rect 111886 343544 111892 343596
rect 111944 343584 111950 343596
rect 119982 343584 119988 343596
rect 111944 343556 119988 343584
rect 111944 343544 111950 343556
rect 119982 343544 119988 343556
rect 120040 343544 120046 343596
rect 115842 342864 115848 342916
rect 115900 342904 115906 342916
rect 277394 342904 277400 342916
rect 115900 342876 277400 342904
rect 115900 342864 115906 342876
rect 277394 342864 277400 342876
rect 277452 342864 277458 342916
rect 111886 342184 111892 342236
rect 111944 342224 111950 342236
rect 117222 342224 117228 342236
rect 111944 342196 117228 342224
rect 111944 342184 111950 342196
rect 117222 342184 117228 342196
rect 117280 342184 117286 342236
rect 124950 341504 124956 341556
rect 125008 341544 125014 341556
rect 580258 341544 580264 341556
rect 125008 341516 580264 341544
rect 125008 341504 125014 341516
rect 580258 341504 580264 341516
rect 580316 341504 580322 341556
rect 65886 340892 65892 340944
rect 65944 340932 65950 340944
rect 67634 340932 67640 340944
rect 65944 340904 67640 340932
rect 65944 340892 65950 340904
rect 67634 340892 67640 340904
rect 67692 340892 67698 340944
rect 117222 340892 117228 340944
rect 117280 340932 117286 340944
rect 120718 340932 120724 340944
rect 117280 340904 120724 340932
rect 117280 340892 117286 340904
rect 120718 340892 120724 340904
rect 120776 340892 120782 340944
rect 110322 340144 110328 340196
rect 110380 340184 110386 340196
rect 112162 340184 112168 340196
rect 110380 340156 112168 340184
rect 110380 340144 110386 340156
rect 112162 340144 112168 340156
rect 112220 340144 112226 340196
rect 395338 340184 395344 340196
rect 113146 340156 395344 340184
rect 70486 339940 70492 339992
rect 70544 339980 70550 339992
rect 79318 339980 79324 339992
rect 70544 339952 79324 339980
rect 70544 339940 70550 339952
rect 79318 339940 79324 339952
rect 79376 339940 79382 339992
rect 107562 339940 107568 339992
rect 107620 339980 107626 339992
rect 113146 339980 113174 340156
rect 395338 340144 395344 340156
rect 395396 340144 395402 340196
rect 107620 339952 113174 339980
rect 107620 339940 107626 339952
rect 4798 339396 4804 339448
rect 4856 339436 4862 339448
rect 83550 339436 83556 339448
rect 4856 339408 83556 339436
rect 4856 339396 4862 339408
rect 83550 339396 83556 339408
rect 83608 339396 83614 339448
rect 84838 339396 84844 339448
rect 84896 339436 84902 339448
rect 316770 339436 316776 339448
rect 84896 339408 316776 339436
rect 84896 339396 84902 339408
rect 316770 339396 316776 339408
rect 316828 339396 316834 339448
rect 65978 339328 65984 339380
rect 66036 339368 66042 339380
rect 125686 339368 125692 339380
rect 66036 339340 125692 339368
rect 66036 339328 66042 339340
rect 125686 339328 125692 339340
rect 125744 339368 125750 339380
rect 126238 339368 126244 339380
rect 125744 339340 126244 339368
rect 125744 339328 125750 339340
rect 126238 339328 126244 339340
rect 126296 339328 126302 339380
rect 58618 339260 58624 339312
rect 58676 339300 58682 339312
rect 91094 339300 91100 339312
rect 58676 339272 91100 339300
rect 58676 339260 58682 339272
rect 91094 339260 91100 339272
rect 91152 339300 91158 339312
rect 91922 339300 91928 339312
rect 91152 339272 91928 339300
rect 91152 339260 91158 339272
rect 91922 339260 91928 339272
rect 91980 339260 91986 339312
rect 95142 339260 95148 339312
rect 95200 339300 95206 339312
rect 117314 339300 117320 339312
rect 95200 339272 117320 339300
rect 95200 339260 95206 339272
rect 117314 339260 117320 339272
rect 117372 339260 117378 339312
rect 106274 338852 106280 338904
rect 106332 338892 106338 338904
rect 109586 338892 109592 338904
rect 106332 338864 109592 338892
rect 106332 338852 106338 338864
rect 109586 338852 109592 338864
rect 109644 338852 109650 338904
rect 105538 338784 105544 338836
rect 105596 338824 105602 338836
rect 113358 338824 113364 338836
rect 105596 338796 113364 338824
rect 105596 338784 105602 338796
rect 113358 338784 113364 338796
rect 113416 338784 113422 338836
rect 68554 338716 68560 338768
rect 68612 338756 68618 338768
rect 284294 338756 284300 338768
rect 68612 338728 284300 338756
rect 68612 338716 68618 338728
rect 284294 338716 284300 338728
rect 284352 338716 284358 338768
rect 32398 338036 32404 338088
rect 32456 338076 32462 338088
rect 98638 338076 98644 338088
rect 32456 338048 98644 338076
rect 32456 338036 32462 338048
rect 98638 338036 98644 338048
rect 98696 338036 98702 338088
rect 104158 338036 104164 338088
rect 104216 338076 104222 338088
rect 115198 338076 115204 338088
rect 104216 338048 115204 338076
rect 104216 338036 104222 338048
rect 115198 338036 115204 338048
rect 115256 338036 115262 338088
rect 129826 338076 129832 338088
rect 122806 338048 129832 338076
rect 66070 337968 66076 338020
rect 66128 338008 66134 338020
rect 73890 338008 73896 338020
rect 66128 337980 73896 338008
rect 66128 337968 66134 337980
rect 73890 337968 73896 337980
rect 73948 337968 73954 338020
rect 78398 337968 78404 338020
rect 78456 338008 78462 338020
rect 122806 338008 122834 338048
rect 129826 338036 129832 338048
rect 129884 338076 129890 338088
rect 130378 338076 130384 338088
rect 129884 338048 130384 338076
rect 129884 338036 129890 338048
rect 130378 338036 130384 338048
rect 130436 338036 130442 338088
rect 78456 337980 122834 338008
rect 78456 337968 78462 337980
rect 80974 337900 80980 337952
rect 81032 337940 81038 337952
rect 107562 337940 107568 337952
rect 81032 337912 107568 337940
rect 81032 337900 81038 337912
rect 107562 337900 107568 337912
rect 107620 337900 107626 337952
rect 84194 337832 84200 337884
rect 84252 337872 84258 337884
rect 90082 337872 90088 337884
rect 84252 337844 90088 337872
rect 84252 337832 84258 337844
rect 90082 337832 90088 337844
rect 90140 337832 90146 337884
rect 70670 337696 70676 337748
rect 70728 337736 70734 337748
rect 72418 337736 72424 337748
rect 70728 337708 72424 337736
rect 70728 337696 70734 337708
rect 72418 337696 72424 337708
rect 72476 337696 72482 337748
rect 100294 337696 100300 337748
rect 100352 337736 100358 337748
rect 101398 337736 101404 337748
rect 100352 337708 101404 337736
rect 100352 337696 100358 337708
rect 101398 337696 101404 337708
rect 101456 337696 101462 337748
rect 71314 337560 71320 337612
rect 71372 337600 71378 337612
rect 73798 337600 73804 337612
rect 71372 337572 73804 337600
rect 71372 337560 71378 337572
rect 73798 337560 73804 337572
rect 73856 337560 73862 337612
rect 87414 337560 87420 337612
rect 87472 337600 87478 337612
rect 89070 337600 89076 337612
rect 87472 337572 89076 337600
rect 87472 337560 87478 337572
rect 89070 337560 89076 337572
rect 89128 337560 89134 337612
rect 100018 337560 100024 337612
rect 100076 337600 100082 337612
rect 114554 337600 114560 337612
rect 100076 337572 114560 337600
rect 100076 337560 100082 337572
rect 114554 337560 114560 337572
rect 114612 337560 114618 337612
rect 109310 337492 109316 337544
rect 109368 337532 109374 337544
rect 191098 337532 191104 337544
rect 109368 337504 191104 337532
rect 109368 337492 109374 337504
rect 191098 337492 191104 337504
rect 191156 337492 191162 337544
rect 73246 337424 73252 337476
rect 73304 337464 73310 337476
rect 80422 337464 80428 337476
rect 73304 337436 80428 337464
rect 73304 337424 73310 337436
rect 80422 337424 80428 337436
rect 80480 337424 80486 337476
rect 81618 337424 81624 337476
rect 81676 337464 81682 337476
rect 188338 337464 188344 337476
rect 81676 337436 188344 337464
rect 81676 337424 81682 337436
rect 188338 337424 188344 337436
rect 188396 337424 188402 337476
rect 74534 337356 74540 337408
rect 74592 337396 74598 337408
rect 87598 337396 87604 337408
rect 74592 337368 87604 337396
rect 74592 337356 74598 337368
rect 87598 337356 87604 337368
rect 87656 337356 87662 337408
rect 92566 337356 92572 337408
rect 92624 337396 92630 337408
rect 307018 337396 307024 337408
rect 92624 337368 307024 337396
rect 92624 337356 92630 337368
rect 307018 337356 307024 337368
rect 307076 337356 307082 337408
rect 70026 336948 70032 337000
rect 70084 336988 70090 337000
rect 75270 336988 75276 337000
rect 70084 336960 75276 336988
rect 70084 336948 70090 336960
rect 75270 336948 75276 336960
rect 75328 336948 75334 337000
rect 72602 336744 72608 336796
rect 72660 336784 72666 336796
rect 75178 336784 75184 336796
rect 72660 336756 75184 336784
rect 72660 336744 72666 336756
rect 75178 336744 75184 336756
rect 75236 336744 75242 336796
rect 35250 336676 35256 336728
rect 35308 336716 35314 336728
rect 95878 336716 95884 336728
rect 35308 336688 95884 336716
rect 35308 336676 35314 336688
rect 95878 336676 95884 336688
rect 95936 336716 95942 336728
rect 96430 336716 96436 336728
rect 95936 336688 96436 336716
rect 95936 336676 95942 336688
rect 96430 336676 96436 336688
rect 96488 336676 96494 336728
rect 68830 336132 68836 336184
rect 68888 336172 68894 336184
rect 269114 336172 269120 336184
rect 68888 336144 269120 336172
rect 68888 336132 68894 336144
rect 269114 336132 269120 336144
rect 269172 336132 269178 336184
rect 60458 336064 60464 336116
rect 60516 336104 60522 336116
rect 88978 336104 88984 336116
rect 60516 336076 88984 336104
rect 60516 336064 60522 336076
rect 88978 336064 88984 336076
rect 89036 336064 89042 336116
rect 90082 336064 90088 336116
rect 90140 336104 90146 336116
rect 343634 336104 343640 336116
rect 90140 336076 343640 336104
rect 90140 336064 90146 336076
rect 343634 336064 343640 336076
rect 343692 336064 343698 336116
rect 88702 335996 88708 336048
rect 88760 336036 88766 336048
rect 126974 336036 126980 336048
rect 88760 336008 126980 336036
rect 88760 335996 88766 336008
rect 126974 335996 126980 336008
rect 127032 336036 127038 336048
rect 582374 336036 582380 336048
rect 127032 336008 582380 336036
rect 127032 335996 127038 336008
rect 582374 335996 582380 336008
rect 582432 335996 582438 336048
rect 56318 334840 56324 334892
rect 56376 334880 56382 334892
rect 82906 334880 82912 334892
rect 56376 334852 82912 334880
rect 56376 334840 56382 334852
rect 82906 334840 82912 334852
rect 82964 334840 82970 334892
rect 57698 334772 57704 334824
rect 57756 334812 57762 334824
rect 94498 334812 94504 334824
rect 57756 334784 94504 334812
rect 57756 334772 57762 334784
rect 94498 334772 94504 334784
rect 94556 334772 94562 334824
rect 99650 334744 99656 334756
rect 55186 334716 99656 334744
rect 3418 334568 3424 334620
rect 3476 334608 3482 334620
rect 53558 334608 53564 334620
rect 3476 334580 53564 334608
rect 3476 334568 3482 334580
rect 53558 334568 53564 334580
rect 53616 334608 53622 334620
rect 55186 334608 55214 334716
rect 99650 334704 99656 334716
rect 99708 334704 99714 334756
rect 99742 334704 99748 334756
rect 99800 334744 99806 334756
rect 112070 334744 112076 334756
rect 99800 334716 112076 334744
rect 99800 334704 99806 334716
rect 112070 334704 112076 334716
rect 112128 334744 112134 334756
rect 131114 334744 131120 334756
rect 112128 334716 131120 334744
rect 112128 334704 112134 334716
rect 131114 334704 131120 334716
rect 131172 334704 131178 334756
rect 61930 334636 61936 334688
rect 61988 334676 61994 334688
rect 133874 334676 133880 334688
rect 61988 334648 133880 334676
rect 61988 334636 61994 334648
rect 133874 334636 133880 334648
rect 133932 334636 133938 334688
rect 53616 334580 55214 334608
rect 53616 334568 53622 334580
rect 68738 334568 68744 334620
rect 68796 334608 68802 334620
rect 309870 334608 309876 334620
rect 68796 334580 309876 334608
rect 68796 334568 68802 334580
rect 309870 334568 309876 334580
rect 309928 334568 309934 334620
rect 107378 333888 107384 333940
rect 107436 333928 107442 333940
rect 341518 333928 341524 333940
rect 107436 333900 341524 333928
rect 107436 333888 107442 333900
rect 341518 333888 341524 333900
rect 341576 333888 341582 333940
rect 25498 333820 25504 333872
rect 25556 333860 25562 333872
rect 107746 333860 107752 333872
rect 25556 333832 107752 333860
rect 25556 333820 25562 333832
rect 107746 333820 107752 333832
rect 107804 333820 107810 333872
rect 67358 333208 67364 333260
rect 67416 333248 67422 333260
rect 273254 333248 273260 333260
rect 67416 333220 273260 333248
rect 67416 333208 67422 333220
rect 273254 333208 273260 333220
rect 273312 333208 273318 333260
rect 106918 332596 106924 332648
rect 106976 332636 106982 332648
rect 107378 332636 107384 332648
rect 106976 332608 107384 332636
rect 106976 332596 106982 332608
rect 107378 332596 107384 332608
rect 107436 332596 107442 332648
rect 39298 332528 39304 332580
rect 39356 332568 39362 332580
rect 99742 332568 99748 332580
rect 39356 332540 99748 332568
rect 39356 332528 39362 332540
rect 99742 332528 99748 332540
rect 99800 332528 99806 332580
rect 52270 331848 52276 331900
rect 52328 331888 52334 331900
rect 91278 331888 91284 331900
rect 52328 331860 91284 331888
rect 52328 331848 52334 331860
rect 91278 331848 91284 331860
rect 91336 331848 91342 331900
rect 80422 331168 80428 331220
rect 80480 331208 80486 331220
rect 124306 331208 124312 331220
rect 80480 331180 124312 331208
rect 80480 331168 80486 331180
rect 124306 331168 124312 331180
rect 124364 331208 124370 331220
rect 124950 331208 124956 331220
rect 124364 331180 124956 331208
rect 124364 331168 124370 331180
rect 124950 331168 124956 331180
rect 125008 331168 125014 331220
rect 61930 330556 61936 330608
rect 61988 330596 61994 330608
rect 113266 330596 113272 330608
rect 61988 330568 113272 330596
rect 61988 330556 61994 330568
rect 113266 330556 113272 330568
rect 113324 330556 113330 330608
rect 98362 330488 98368 330540
rect 98420 330528 98426 330540
rect 293954 330528 293960 330540
rect 98420 330500 293960 330528
rect 98420 330488 98426 330500
rect 293954 330488 293960 330500
rect 294012 330488 294018 330540
rect 67450 329196 67456 329248
rect 67508 329236 67514 329248
rect 115198 329236 115204 329248
rect 67508 329208 115204 329236
rect 67508 329196 67514 329208
rect 115198 329196 115204 329208
rect 115256 329196 115262 329248
rect 39850 329128 39856 329180
rect 39908 329168 39914 329180
rect 102870 329168 102876 329180
rect 39908 329140 102876 329168
rect 39908 329128 39914 329140
rect 102870 329128 102876 329140
rect 102928 329128 102934 329180
rect 69106 329060 69112 329112
rect 69164 329100 69170 329112
rect 281534 329100 281540 329112
rect 69164 329072 281540 329100
rect 69164 329060 69170 329072
rect 281534 329060 281540 329072
rect 281592 329060 281598 329112
rect 65886 328380 65892 328432
rect 65944 328420 65950 328432
rect 140866 328420 140872 328432
rect 65944 328392 140872 328420
rect 65944 328380 65950 328392
rect 140866 328380 140872 328392
rect 140924 328420 140930 328432
rect 141418 328420 141424 328432
rect 140924 328392 141424 328420
rect 140924 328380 140930 328392
rect 141418 328380 141424 328392
rect 141476 328380 141482 328432
rect 73154 327768 73160 327820
rect 73212 327808 73218 327820
rect 109126 327808 109132 327820
rect 73212 327780 109132 327808
rect 73212 327768 73218 327780
rect 109126 327768 109132 327780
rect 109184 327768 109190 327820
rect 79042 327700 79048 327752
rect 79100 327740 79106 327752
rect 204898 327740 204904 327752
rect 79100 327712 204904 327740
rect 79100 327700 79106 327712
rect 204898 327700 204904 327712
rect 204956 327700 204962 327752
rect 106734 326340 106740 326392
rect 106792 326380 106798 326392
rect 152458 326380 152464 326392
rect 106792 326352 152464 326380
rect 106792 326340 106798 326352
rect 152458 326340 152464 326352
rect 152516 326340 152522 326392
rect 73890 324912 73896 324964
rect 73948 324952 73954 324964
rect 114554 324952 114560 324964
rect 73948 324924 114560 324952
rect 73948 324912 73954 324924
rect 114554 324912 114560 324924
rect 114612 324912 114618 324964
rect 102134 323688 102140 323740
rect 102192 323728 102198 323740
rect 121546 323728 121552 323740
rect 102192 323700 121552 323728
rect 102192 323688 102198 323700
rect 121546 323688 121552 323700
rect 121604 323728 121610 323740
rect 121822 323728 121828 323740
rect 121604 323700 121828 323728
rect 121604 323688 121610 323700
rect 121822 323688 121828 323700
rect 121880 323688 121886 323740
rect 97074 323620 97080 323672
rect 97132 323660 97138 323672
rect 284386 323660 284392 323672
rect 97132 323632 284392 323660
rect 97132 323620 97138 323632
rect 284386 323620 284392 323632
rect 284444 323620 284450 323672
rect 84286 323552 84292 323604
rect 84344 323592 84350 323604
rect 109494 323592 109500 323604
rect 84344 323564 109500 323592
rect 84344 323552 84350 323564
rect 109494 323552 109500 323564
rect 109552 323552 109558 323604
rect 121822 323552 121828 323604
rect 121880 323592 121886 323604
rect 582558 323592 582564 323604
rect 121880 323564 582564 323592
rect 121880 323552 121886 323564
rect 582558 323552 582564 323564
rect 582616 323552 582622 323604
rect 71038 322328 71044 322380
rect 71096 322368 71102 322380
rect 102134 322368 102140 322380
rect 71096 322340 102140 322368
rect 71096 322328 71102 322340
rect 102134 322328 102140 322340
rect 102192 322328 102198 322380
rect 93854 322260 93860 322312
rect 93912 322300 93918 322312
rect 287054 322300 287060 322312
rect 93912 322272 287060 322300
rect 93912 322260 93918 322272
rect 287054 322260 287060 322272
rect 287112 322260 287118 322312
rect 68922 322192 68928 322244
rect 68980 322232 68986 322244
rect 308398 322232 308404 322244
rect 68980 322204 308404 322232
rect 68980 322192 68986 322204
rect 308398 322192 308404 322204
rect 308456 322192 308462 322244
rect 101398 320832 101404 320884
rect 101456 320872 101462 320884
rect 349246 320872 349252 320884
rect 101456 320844 349252 320872
rect 101456 320832 101462 320844
rect 349246 320832 349252 320844
rect 349304 320832 349310 320884
rect 79318 319472 79324 319524
rect 79376 319512 79382 319524
rect 155218 319512 155224 319524
rect 79376 319484 155224 319512
rect 79376 319472 79382 319484
rect 155218 319472 155224 319484
rect 155276 319472 155282 319524
rect 59170 319404 59176 319456
rect 59228 319444 59234 319456
rect 197998 319444 198004 319456
rect 59228 319416 198004 319444
rect 59228 319404 59234 319416
rect 197998 319404 198004 319416
rect 198056 319404 198062 319456
rect 95142 318724 95148 318776
rect 95200 318764 95206 318776
rect 101398 318764 101404 318776
rect 95200 318736 101404 318764
rect 95200 318724 95206 318736
rect 101398 318724 101404 318736
rect 101456 318724 101462 318776
rect 77110 318044 77116 318096
rect 77168 318084 77174 318096
rect 204990 318084 204996 318096
rect 77168 318056 204996 318084
rect 77168 318044 77174 318056
rect 204990 318044 204996 318056
rect 205048 318044 205054 318096
rect 128998 317364 129004 317416
rect 129056 317404 129062 317416
rect 131206 317404 131212 317416
rect 129056 317376 131212 317404
rect 129056 317364 129062 317376
rect 131206 317364 131212 317376
rect 131264 317404 131270 317416
rect 580166 317404 580172 317416
rect 131264 317376 580172 317404
rect 131264 317364 131270 317376
rect 580166 317364 580172 317376
rect 580224 317364 580230 317416
rect 64598 316820 64604 316872
rect 64656 316860 64662 316872
rect 124398 316860 124404 316872
rect 64656 316832 124404 316860
rect 64656 316820 64662 316832
rect 124398 316820 124404 316832
rect 124456 316820 124462 316872
rect 61838 316752 61844 316804
rect 61896 316792 61902 316804
rect 134058 316792 134064 316804
rect 61896 316764 134064 316792
rect 61896 316752 61902 316764
rect 134058 316752 134064 316764
rect 134116 316752 134122 316804
rect 76466 316684 76472 316736
rect 76524 316724 76530 316736
rect 213178 316724 213184 316736
rect 76524 316696 213184 316724
rect 76524 316684 76530 316696
rect 213178 316684 213184 316696
rect 213236 316684 213242 316736
rect 89346 315256 89352 315308
rect 89404 315296 89410 315308
rect 146938 315296 146944 315308
rect 89404 315268 146944 315296
rect 89404 315256 89410 315268
rect 146938 315256 146944 315268
rect 146996 315256 147002 315308
rect 63126 314032 63132 314084
rect 63184 314072 63190 314084
rect 84838 314072 84844 314084
rect 63184 314044 84844 314072
rect 63184 314032 63190 314044
rect 84838 314032 84844 314044
rect 84896 314032 84902 314084
rect 94498 313964 94504 314016
rect 94556 314004 94562 314016
rect 108666 314004 108672 314016
rect 94556 313976 108672 314004
rect 94556 313964 94562 313976
rect 108666 313964 108672 313976
rect 108724 313964 108730 314016
rect 63402 313896 63408 313948
rect 63460 313936 63466 313948
rect 129918 313936 129924 313948
rect 63460 313908 129924 313936
rect 63460 313896 63466 313908
rect 129918 313896 129924 313908
rect 129976 313896 129982 313948
rect 71958 312604 71964 312656
rect 72016 312644 72022 312656
rect 287698 312644 287704 312656
rect 72016 312616 287704 312644
rect 72016 312604 72022 312616
rect 287698 312604 287704 312616
rect 287756 312604 287762 312656
rect 3418 312536 3424 312588
rect 3476 312576 3482 312588
rect 115934 312576 115940 312588
rect 3476 312548 115940 312576
rect 3476 312536 3482 312548
rect 115934 312536 115940 312548
rect 115992 312536 115998 312588
rect 580166 312576 580172 312588
rect 132466 312548 580172 312576
rect 124398 312468 124404 312520
rect 124456 312508 124462 312520
rect 124858 312508 124864 312520
rect 124456 312480 124864 312508
rect 124456 312468 124462 312480
rect 124858 312468 124864 312480
rect 124916 312508 124922 312520
rect 132466 312508 132494 312548
rect 580166 312536 580172 312548
rect 580224 312536 580230 312588
rect 124916 312480 132494 312508
rect 124916 312468 124922 312480
rect 72418 311176 72424 311228
rect 72476 311216 72482 311228
rect 103514 311216 103520 311228
rect 72476 311188 103520 311216
rect 72476 311176 72482 311188
rect 103514 311176 103520 311188
rect 103572 311176 103578 311228
rect 79686 311108 79692 311160
rect 79744 311148 79750 311160
rect 180058 311148 180064 311160
rect 79744 311120 180064 311148
rect 79744 311108 79750 311120
rect 180058 311108 180064 311120
rect 180116 311108 180122 311160
rect 75914 310496 75920 310548
rect 75972 310536 75978 310548
rect 295978 310536 295984 310548
rect 75972 310508 295984 310536
rect 75972 310496 75978 310508
rect 295978 310496 295984 310508
rect 296036 310496 296042 310548
rect 75822 309816 75828 309868
rect 75880 309856 75886 309868
rect 121638 309856 121644 309868
rect 75880 309828 121644 309856
rect 75880 309816 75886 309828
rect 121638 309816 121644 309828
rect 121696 309816 121702 309868
rect 75270 309748 75276 309800
rect 75328 309788 75334 309800
rect 291194 309788 291200 309800
rect 75328 309760 291200 309788
rect 75328 309748 75334 309760
rect 291194 309748 291200 309760
rect 291252 309748 291258 309800
rect 101582 308660 101588 308712
rect 101640 308700 101646 308712
rect 113818 308700 113824 308712
rect 101640 308672 113824 308700
rect 101640 308660 101646 308672
rect 113818 308660 113824 308672
rect 113876 308660 113882 308712
rect 87598 308592 87604 308644
rect 87656 308632 87662 308644
rect 106918 308632 106924 308644
rect 87656 308604 106924 308632
rect 87656 308592 87662 308604
rect 106918 308592 106924 308604
rect 106976 308592 106982 308644
rect 89070 308524 89076 308576
rect 89128 308564 89134 308576
rect 274634 308564 274640 308576
rect 89128 308536 274640 308564
rect 89128 308524 89134 308536
rect 274634 308524 274640 308536
rect 274692 308524 274698 308576
rect 69014 308456 69020 308508
rect 69072 308496 69078 308508
rect 298094 308496 298100 308508
rect 69072 308468 298100 308496
rect 69072 308456 69078 308468
rect 298094 308456 298100 308468
rect 298152 308456 298158 308508
rect 80054 308388 80060 308440
rect 80112 308428 80118 308440
rect 121454 308428 121460 308440
rect 80112 308400 121460 308428
rect 80112 308388 80118 308400
rect 121454 308388 121460 308400
rect 121512 308428 121518 308440
rect 582834 308428 582840 308440
rect 121512 308400 582840 308428
rect 121512 308388 121518 308400
rect 582834 308388 582840 308400
rect 582892 308388 582898 308440
rect 76558 307096 76564 307148
rect 76616 307136 76622 307148
rect 159358 307136 159364 307148
rect 76616 307108 159364 307136
rect 76616 307096 76622 307108
rect 159358 307096 159364 307108
rect 159416 307096 159422 307148
rect 88058 307028 88064 307080
rect 88116 307068 88122 307080
rect 278774 307068 278780 307080
rect 88116 307040 278780 307068
rect 88116 307028 88122 307040
rect 278774 307028 278780 307040
rect 278832 307028 278838 307080
rect 81434 306416 81440 306468
rect 81492 306456 81498 306468
rect 246298 306456 246304 306468
rect 81492 306428 246304 306456
rect 81492 306416 81498 306428
rect 246298 306416 246304 306428
rect 246356 306416 246362 306468
rect 89714 306348 89720 306400
rect 89772 306388 89778 306400
rect 300118 306388 300124 306400
rect 89772 306360 300124 306388
rect 89772 306348 89778 306360
rect 300118 306348 300124 306360
rect 300176 306348 300182 306400
rect 3418 306280 3424 306332
rect 3476 306320 3482 306332
rect 42702 306320 42708 306332
rect 3476 306292 42708 306320
rect 3476 306280 3482 306292
rect 42702 306280 42708 306292
rect 42760 306280 42766 306332
rect 95878 305804 95884 305856
rect 95936 305844 95942 305856
rect 123110 305844 123116 305856
rect 95936 305816 123116 305844
rect 95936 305804 95942 305816
rect 123110 305804 123116 305816
rect 123168 305804 123174 305856
rect 61838 305736 61844 305788
rect 61896 305776 61902 305788
rect 110414 305776 110420 305788
rect 61896 305748 110420 305776
rect 61896 305736 61902 305748
rect 110414 305736 110420 305748
rect 110472 305736 110478 305788
rect 42702 305668 42708 305720
rect 42760 305708 42766 305720
rect 117406 305708 117412 305720
rect 42760 305680 117412 305708
rect 42760 305668 42766 305680
rect 117406 305668 117412 305680
rect 117464 305668 117470 305720
rect 86126 305600 86132 305652
rect 86184 305640 86190 305652
rect 217318 305640 217324 305652
rect 86184 305612 217324 305640
rect 86184 305600 86190 305612
rect 217318 305600 217324 305612
rect 217376 305600 217382 305652
rect 88334 304988 88340 305040
rect 88392 305028 88398 305040
rect 356054 305028 356060 305040
rect 88392 305000 356060 305028
rect 88392 304988 88398 305000
rect 356054 304988 356060 305000
rect 356112 304988 356118 305040
rect 72234 304240 72240 304292
rect 72292 304280 72298 304292
rect 124214 304280 124220 304292
rect 72292 304252 124220 304280
rect 72292 304240 72298 304252
rect 124214 304240 124220 304252
rect 124272 304240 124278 304292
rect 106090 303764 106096 303816
rect 106148 303804 106154 303816
rect 110506 303804 110512 303816
rect 106148 303776 110512 303804
rect 106148 303764 106154 303776
rect 110506 303764 110512 303776
rect 110564 303764 110570 303816
rect 111702 303764 111708 303816
rect 111760 303804 111766 303816
rect 111886 303804 111892 303816
rect 111760 303776 111892 303804
rect 111760 303764 111766 303776
rect 111886 303764 111892 303776
rect 111944 303764 111950 303816
rect 116670 303764 116676 303816
rect 116728 303804 116734 303816
rect 117314 303804 117320 303816
rect 116728 303776 117320 303804
rect 116728 303764 116734 303776
rect 117314 303764 117320 303776
rect 117372 303764 117378 303816
rect 79318 303696 79324 303748
rect 79376 303736 79382 303748
rect 229738 303736 229744 303748
rect 79376 303708 229744 303736
rect 79376 303696 79382 303708
rect 229738 303696 229744 303708
rect 229796 303696 229802 303748
rect 67450 303628 67456 303680
rect 67508 303668 67514 303680
rect 226978 303668 226984 303680
rect 67508 303640 226984 303668
rect 67508 303628 67514 303640
rect 226978 303628 226984 303640
rect 227036 303628 227042 303680
rect 69014 302948 69020 303000
rect 69072 302988 69078 303000
rect 111794 302988 111800 303000
rect 69072 302960 111800 302988
rect 69072 302948 69078 302960
rect 111794 302948 111800 302960
rect 111852 302948 111858 303000
rect 86770 302880 86776 302932
rect 86828 302920 86834 302932
rect 151078 302920 151084 302932
rect 86828 302892 151084 302920
rect 86828 302880 86834 302892
rect 151078 302880 151084 302892
rect 151136 302880 151142 302932
rect 100846 302404 100852 302456
rect 100904 302444 100910 302456
rect 244918 302444 244924 302456
rect 100904 302416 244924 302444
rect 100904 302404 100910 302416
rect 244918 302404 244924 302416
rect 244976 302404 244982 302456
rect 74534 302336 74540 302388
rect 74592 302376 74598 302388
rect 222838 302376 222844 302388
rect 74592 302348 222844 302376
rect 74592 302336 74598 302348
rect 222838 302336 222844 302348
rect 222896 302336 222902 302388
rect 106366 302268 106372 302320
rect 106424 302308 106430 302320
rect 319438 302308 319444 302320
rect 106424 302280 319444 302308
rect 106424 302268 106430 302280
rect 319438 302268 319444 302280
rect 319496 302268 319502 302320
rect 103606 302200 103612 302252
rect 103664 302240 103670 302252
rect 349338 302240 349344 302252
rect 103664 302212 349344 302240
rect 103664 302200 103670 302212
rect 349338 302200 349344 302212
rect 349396 302200 349402 302252
rect 122098 302132 122104 302184
rect 122156 302172 122162 302184
rect 124214 302172 124220 302184
rect 122156 302144 124220 302172
rect 122156 302132 122162 302144
rect 124214 302132 124220 302144
rect 124272 302132 124278 302184
rect 66070 301452 66076 301504
rect 66128 301492 66134 301504
rect 111702 301492 111708 301504
rect 66128 301464 111708 301492
rect 66128 301452 66134 301464
rect 111702 301452 111708 301464
rect 111760 301492 111766 301504
rect 583110 301492 583116 301504
rect 111760 301464 583116 301492
rect 111760 301452 111766 301464
rect 583110 301452 583116 301464
rect 583168 301452 583174 301504
rect 102134 300976 102140 301028
rect 102192 301016 102198 301028
rect 199378 301016 199384 301028
rect 102192 300988 199384 301016
rect 102192 300976 102198 300988
rect 199378 300976 199384 300988
rect 199436 300976 199442 301028
rect 73246 300908 73252 300960
rect 73304 300948 73310 300960
rect 192478 300948 192484 300960
rect 73304 300920 192484 300948
rect 73304 300908 73310 300920
rect 192478 300908 192484 300920
rect 192536 300908 192542 300960
rect 85574 300840 85580 300892
rect 85632 300880 85638 300892
rect 224218 300880 224224 300892
rect 85632 300852 224224 300880
rect 85632 300840 85638 300852
rect 224218 300840 224224 300852
rect 224276 300840 224282 300892
rect 52178 300160 52184 300212
rect 52236 300200 52242 300212
rect 97994 300200 98000 300212
rect 52236 300172 98000 300200
rect 52236 300160 52242 300172
rect 97994 300160 98000 300172
rect 98052 300160 98058 300212
rect 63310 300092 63316 300144
rect 63368 300132 63374 300144
rect 132678 300132 132684 300144
rect 63368 300104 132684 300132
rect 63368 300092 63374 300104
rect 132678 300092 132684 300104
rect 132736 300092 132742 300144
rect 102318 299752 102324 299804
rect 102376 299792 102382 299804
rect 213270 299792 213276 299804
rect 102376 299764 213276 299792
rect 102376 299752 102382 299764
rect 213270 299752 213276 299764
rect 213328 299752 213334 299804
rect 89806 299684 89812 299736
rect 89864 299724 89870 299736
rect 232590 299724 232596 299736
rect 89864 299696 232596 299724
rect 89864 299684 89870 299696
rect 232590 299684 232596 299696
rect 232648 299684 232654 299736
rect 80606 299616 80612 299668
rect 80664 299656 80670 299668
rect 238018 299656 238024 299668
rect 80664 299628 238024 299656
rect 80664 299616 80670 299628
rect 238018 299616 238024 299628
rect 238076 299616 238082 299668
rect 97350 299548 97356 299600
rect 97408 299588 97414 299600
rect 333238 299588 333244 299600
rect 97408 299560 333244 299588
rect 97408 299548 97414 299560
rect 333238 299548 333244 299560
rect 333296 299548 333302 299600
rect 88426 299480 88432 299532
rect 88484 299520 88490 299532
rect 335354 299520 335360 299532
rect 88484 299492 335360 299520
rect 88484 299480 88490 299492
rect 335354 299480 335360 299492
rect 335412 299480 335418 299532
rect 83458 298800 83464 298852
rect 83516 298840 83522 298852
rect 127158 298840 127164 298852
rect 83516 298812 127164 298840
rect 83516 298800 83522 298812
rect 127158 298800 127164 298812
rect 127216 298800 127222 298852
rect 60458 298732 60464 298784
rect 60516 298772 60522 298784
rect 105538 298772 105544 298784
rect 60516 298744 105544 298772
rect 60516 298732 60522 298744
rect 105538 298732 105544 298744
rect 105596 298732 105602 298784
rect 84194 298392 84200 298444
rect 84252 298432 84258 298444
rect 144178 298432 144184 298444
rect 84252 298404 144184 298432
rect 84252 298392 84258 298404
rect 144178 298392 144184 298404
rect 144236 298392 144242 298444
rect 87414 298324 87420 298376
rect 87472 298364 87478 298376
rect 210510 298364 210516 298376
rect 87472 298336 210516 298364
rect 87472 298324 87478 298336
rect 210510 298324 210516 298336
rect 210568 298324 210574 298376
rect 111242 298256 111248 298308
rect 111300 298296 111306 298308
rect 318058 298296 318064 298308
rect 111300 298268 318064 298296
rect 111300 298256 111306 298268
rect 318058 298256 318064 298268
rect 318116 298256 318122 298308
rect 111886 298188 111892 298240
rect 111944 298228 111950 298240
rect 343726 298228 343732 298240
rect 111944 298200 343732 298228
rect 111944 298188 111950 298200
rect 343726 298188 343732 298200
rect 343784 298188 343790 298240
rect 86770 298120 86776 298172
rect 86828 298160 86834 298172
rect 320818 298160 320824 298172
rect 86828 298132 320824 298160
rect 86828 298120 86834 298132
rect 320818 298120 320824 298132
rect 320876 298120 320882 298172
rect 117406 298052 117412 298104
rect 117464 298092 117470 298104
rect 121546 298092 121552 298104
rect 117464 298064 121552 298092
rect 117464 298052 117470 298064
rect 121546 298052 121552 298064
rect 121604 298052 121610 298104
rect 94498 297440 94504 297492
rect 94556 297480 94562 297492
rect 107746 297480 107752 297492
rect 94556 297452 107752 297480
rect 94556 297440 94562 297452
rect 107746 297440 107752 297452
rect 107804 297440 107810 297492
rect 98638 297372 98644 297424
rect 98696 297412 98702 297424
rect 125870 297412 125876 297424
rect 98696 297384 125876 297412
rect 98696 297372 98702 297384
rect 125870 297372 125876 297384
rect 125928 297372 125934 297424
rect 112530 296896 112536 296948
rect 112588 296936 112594 296948
rect 202230 296936 202236 296948
rect 112588 296908 202236 296936
rect 112588 296896 112594 296908
rect 202230 296896 202236 296908
rect 202288 296896 202294 296948
rect 67542 296828 67548 296880
rect 67600 296868 67606 296880
rect 207658 296868 207664 296880
rect 67600 296840 207664 296868
rect 67600 296828 67606 296840
rect 207658 296828 207664 296840
rect 207716 296828 207722 296880
rect 3418 296760 3424 296812
rect 3476 296800 3482 296812
rect 100018 296800 100024 296812
rect 3476 296772 100024 296800
rect 3476 296760 3482 296772
rect 100018 296760 100024 296772
rect 100076 296760 100082 296812
rect 108666 296760 108672 296812
rect 108724 296800 108730 296812
rect 114646 296800 114652 296812
rect 108724 296772 114652 296800
rect 108724 296760 108730 296772
rect 114646 296760 114652 296772
rect 114704 296760 114710 296812
rect 117038 296760 117044 296812
rect 117096 296800 117102 296812
rect 342346 296800 342352 296812
rect 117096 296772 342352 296800
rect 117096 296760 117102 296772
rect 342346 296760 342352 296772
rect 342404 296760 342410 296812
rect 99006 296692 99012 296744
rect 99064 296732 99070 296744
rect 358814 296732 358820 296744
rect 99064 296704 358820 296732
rect 99064 296692 99070 296704
rect 358814 296692 358820 296704
rect 358872 296692 358878 296744
rect 11698 295944 11704 295996
rect 11756 295984 11762 295996
rect 71314 295984 71320 295996
rect 11756 295956 71320 295984
rect 11756 295944 11762 295956
rect 71314 295944 71320 295956
rect 71372 295984 71378 295996
rect 72418 295984 72424 295996
rect 71372 295956 72424 295984
rect 71372 295944 71378 295956
rect 72418 295944 72424 295956
rect 72476 295944 72482 295996
rect 82906 295672 82912 295724
rect 82964 295712 82970 295724
rect 141418 295712 141424 295724
rect 82964 295684 141424 295712
rect 82964 295672 82970 295684
rect 141418 295672 141424 295684
rect 141476 295672 141482 295724
rect 40678 295604 40684 295656
rect 40736 295644 40742 295656
rect 117314 295644 117320 295656
rect 40736 295616 117320 295644
rect 40736 295604 40742 295616
rect 117314 295604 117320 295616
rect 117372 295644 117378 295656
rect 118326 295644 118332 295656
rect 117372 295616 118332 295644
rect 117372 295604 117378 295616
rect 118326 295604 118332 295616
rect 118384 295604 118390 295656
rect 93210 295536 93216 295588
rect 93268 295576 93274 295588
rect 203518 295576 203524 295588
rect 93268 295548 203524 295576
rect 93268 295536 93274 295548
rect 203518 295536 203524 295548
rect 203576 295536 203582 295588
rect 83550 295468 83556 295520
rect 83608 295508 83614 295520
rect 247678 295508 247684 295520
rect 83608 295480 247684 295508
rect 83608 295468 83614 295480
rect 247678 295468 247684 295480
rect 247736 295468 247742 295520
rect 65978 295400 65984 295452
rect 66036 295440 66042 295452
rect 240778 295440 240784 295452
rect 66036 295412 240784 295440
rect 66036 295400 66042 295412
rect 240778 295400 240784 295412
rect 240836 295400 240842 295452
rect 109310 295332 109316 295384
rect 109368 295372 109374 295384
rect 319530 295372 319536 295384
rect 109368 295344 319536 295372
rect 109368 295332 109374 295344
rect 319530 295332 319536 295344
rect 319588 295332 319594 295384
rect 101398 295264 101404 295316
rect 101456 295304 101462 295316
rect 104802 295304 104808 295316
rect 101456 295276 104808 295304
rect 101456 295264 101462 295276
rect 104802 295264 104808 295276
rect 104860 295264 104866 295316
rect 92750 295128 92756 295180
rect 92808 295168 92814 295180
rect 94406 295168 94412 295180
rect 92808 295140 94412 295168
rect 92808 295128 92814 295140
rect 94406 295128 94412 295140
rect 94464 295128 94470 295180
rect 85482 294924 85488 294976
rect 85540 294964 85546 294976
rect 87598 294964 87604 294976
rect 85540 294936 87604 294964
rect 85540 294924 85546 294936
rect 87598 294924 87604 294936
rect 87656 294924 87662 294976
rect 66162 294720 66168 294772
rect 66220 294760 66226 294772
rect 78398 294760 78404 294772
rect 66220 294732 78404 294760
rect 66220 294720 66226 294732
rect 78398 294720 78404 294732
rect 78456 294720 78462 294772
rect 79042 294692 79048 294704
rect 55186 294664 79048 294692
rect 14458 294584 14464 294636
rect 14516 294624 14522 294636
rect 53650 294624 53656 294636
rect 14516 294596 53656 294624
rect 14516 294584 14522 294596
rect 53650 294584 53656 294596
rect 53708 294624 53714 294636
rect 55186 294624 55214 294664
rect 79042 294652 79048 294664
rect 79100 294652 79106 294704
rect 53708 294596 55214 294624
rect 53708 294584 53714 294596
rect 62022 294584 62028 294636
rect 62080 294624 62086 294636
rect 91278 294624 91284 294636
rect 62080 294596 91284 294624
rect 62080 294584 62086 294596
rect 91278 294584 91284 294596
rect 91336 294584 91342 294636
rect 70026 294380 70032 294432
rect 70084 294420 70090 294432
rect 117958 294420 117964 294432
rect 70084 294392 117964 294420
rect 70084 294380 70090 294392
rect 117958 294380 117964 294392
rect 118016 294380 118022 294432
rect 73154 294312 73160 294364
rect 73212 294352 73218 294364
rect 73614 294352 73620 294364
rect 73212 294324 73620 294352
rect 73212 294312 73218 294324
rect 73614 294312 73620 294324
rect 73672 294312 73678 294364
rect 88334 294312 88340 294364
rect 88392 294352 88398 294364
rect 89070 294352 89076 294364
rect 88392 294324 89076 294352
rect 88392 294312 88398 294324
rect 89070 294312 89076 294324
rect 89128 294312 89134 294364
rect 93946 294312 93952 294364
rect 94004 294352 94010 294364
rect 94774 294352 94780 294364
rect 94004 294324 94780 294352
rect 94004 294312 94010 294324
rect 94774 294312 94780 294324
rect 94832 294312 94838 294364
rect 100018 294312 100024 294364
rect 100076 294352 100082 294364
rect 101582 294352 101588 294364
rect 100076 294324 101588 294352
rect 100076 294312 100082 294324
rect 101582 294312 101588 294324
rect 101640 294312 101646 294364
rect 106274 294312 106280 294364
rect 106332 294352 106338 294364
rect 107102 294352 107108 294364
rect 106332 294324 107108 294352
rect 106332 294312 106338 294324
rect 107102 294312 107108 294324
rect 107160 294312 107166 294364
rect 110322 294312 110328 294364
rect 110380 294352 110386 294364
rect 119798 294352 119804 294364
rect 110380 294324 119804 294352
rect 110380 294312 110386 294324
rect 119798 294312 119804 294324
rect 119856 294312 119862 294364
rect 88058 294244 88064 294296
rect 88116 294284 88122 294296
rect 88116 294256 103514 294284
rect 88116 294244 88122 294256
rect 96430 294216 96436 294228
rect 84166 294188 96436 294216
rect 57882 294108 57888 294160
rect 57940 294148 57946 294160
rect 84166 294148 84194 294188
rect 96430 294176 96436 294188
rect 96488 294176 96494 294228
rect 103486 294216 103514 294256
rect 105446 294244 105452 294296
rect 105504 294284 105510 294296
rect 106090 294284 106096 294296
rect 105504 294256 106096 294284
rect 105504 294244 105510 294256
rect 106090 294244 106096 294256
rect 106148 294284 106154 294296
rect 125042 294284 125048 294296
rect 106148 294256 125048 294284
rect 106148 294244 106154 294256
rect 125042 294244 125048 294256
rect 125100 294244 125106 294296
rect 114462 294216 114468 294228
rect 103486 294188 114468 294216
rect 114462 294176 114468 294188
rect 114520 294176 114526 294228
rect 118970 294176 118976 294228
rect 119028 294216 119034 294228
rect 218698 294216 218704 294228
rect 119028 294188 218704 294216
rect 119028 294176 119034 294188
rect 218698 294176 218704 294188
rect 218756 294176 218762 294228
rect 57940 294120 84194 294148
rect 57940 294108 57946 294120
rect 95786 294108 95792 294160
rect 95844 294148 95850 294160
rect 195330 294148 195336 294160
rect 95844 294120 195336 294148
rect 95844 294108 95850 294120
rect 195330 294108 195336 294120
rect 195388 294108 195394 294160
rect 91922 294040 91928 294092
rect 91980 294080 91986 294092
rect 262214 294080 262220 294092
rect 91980 294052 262220 294080
rect 91980 294040 91986 294052
rect 262214 294040 262220 294052
rect 262272 294040 262278 294092
rect 80146 293972 80152 294024
rect 80204 294012 80210 294024
rect 92750 294012 92756 294024
rect 80204 293984 92756 294012
rect 80204 293972 80210 293984
rect 92750 293972 92756 293984
rect 92808 293972 92814 294024
rect 114370 293972 114376 294024
rect 114428 294012 114434 294024
rect 357434 294012 357440 294024
rect 114428 293984 357440 294012
rect 114428 293972 114434 293984
rect 357434 293972 357440 293984
rect 357492 293972 357498 294024
rect 53098 293292 53104 293344
rect 53156 293332 53162 293344
rect 56410 293332 56416 293344
rect 53156 293304 56416 293332
rect 53156 293292 53162 293304
rect 56410 293292 56416 293304
rect 56468 293332 56474 293344
rect 97074 293332 97080 293344
rect 56468 293304 97080 293332
rect 56468 293292 56474 293304
rect 97074 293292 97080 293304
rect 97132 293292 97138 293344
rect 3602 293224 3608 293276
rect 3660 293264 3666 293276
rect 80146 293264 80152 293276
rect 3660 293236 80152 293264
rect 3660 293224 3666 293236
rect 80146 293224 80152 293236
rect 80204 293224 80210 293276
rect 114462 293224 114468 293276
rect 114520 293264 114526 293276
rect 142798 293264 142804 293276
rect 114520 293236 142804 293264
rect 114520 293224 114526 293236
rect 142798 293224 142804 293236
rect 142856 293224 142862 293276
rect 110598 292816 110604 292868
rect 110656 292856 110662 292868
rect 209222 292856 209228 292868
rect 110656 292828 209228 292856
rect 110656 292816 110662 292828
rect 209222 292816 209228 292828
rect 209280 292816 209286 292868
rect 117682 292748 117688 292800
rect 117740 292788 117746 292800
rect 216122 292788 216128 292800
rect 117740 292760 216128 292788
rect 117740 292748 117746 292760
rect 216122 292748 216128 292760
rect 216180 292748 216186 292800
rect 93854 292680 93860 292732
rect 93912 292720 93918 292732
rect 231118 292720 231124 292732
rect 93912 292692 231124 292720
rect 93912 292680 93918 292692
rect 231118 292680 231124 292692
rect 231176 292680 231182 292732
rect 99650 292612 99656 292664
rect 99708 292652 99714 292664
rect 276106 292652 276112 292664
rect 99708 292624 276112 292652
rect 99708 292612 99714 292624
rect 276106 292612 276112 292624
rect 276164 292612 276170 292664
rect 3510 292544 3516 292596
rect 3568 292584 3574 292596
rect 11698 292584 11704 292596
rect 3568 292556 11704 292584
rect 3568 292544 3574 292556
rect 11698 292544 11704 292556
rect 11756 292544 11762 292596
rect 68646 292544 68652 292596
rect 68704 292584 68710 292596
rect 351914 292584 351920 292596
rect 68704 292556 351920 292584
rect 68704 292544 68710 292556
rect 351914 292544 351920 292556
rect 351972 292544 351978 292596
rect 121454 292476 121460 292528
rect 121512 292516 121518 292528
rect 125594 292516 125600 292528
rect 121512 292488 125600 292516
rect 121512 292476 121518 292488
rect 125594 292476 125600 292488
rect 125652 292476 125658 292528
rect 103514 292068 103520 292120
rect 103572 292068 103578 292120
rect 103532 291224 103560 292068
rect 108298 291864 108304 291916
rect 108356 291904 108362 291916
rect 108356 291876 113174 291904
rect 108356 291864 108362 291876
rect 113146 291292 113174 291876
rect 117958 291864 117964 291916
rect 118016 291904 118022 291916
rect 118016 291876 122834 291904
rect 118016 291864 118022 291876
rect 122806 291836 122834 291876
rect 249058 291836 249064 291848
rect 122806 291808 249064 291836
rect 249058 291796 249064 291808
rect 249116 291796 249122 291848
rect 249150 291292 249156 291304
rect 113146 291264 249156 291292
rect 249150 291252 249156 291264
rect 249208 291252 249214 291304
rect 350626 291224 350632 291236
rect 103532 291196 350632 291224
rect 350626 291184 350632 291196
rect 350684 291184 350690 291236
rect 269758 291116 269764 291168
rect 269816 291156 269822 291168
rect 276014 291156 276020 291168
rect 269816 291128 276020 291156
rect 269816 291116 269822 291128
rect 276014 291116 276020 291128
rect 276072 291116 276078 291168
rect 121454 289892 121460 289944
rect 121512 289932 121518 289944
rect 222930 289932 222936 289944
rect 121512 289904 222936 289932
rect 121512 289892 121518 289904
rect 222930 289892 222936 289904
rect 222988 289892 222994 289944
rect 21358 289824 21364 289876
rect 21416 289864 21422 289876
rect 68002 289864 68008 289876
rect 21416 289836 68008 289864
rect 21416 289824 21422 289836
rect 68002 289824 68008 289836
rect 68060 289824 68066 289876
rect 121730 289824 121736 289876
rect 121788 289864 121794 289876
rect 251818 289864 251824 289876
rect 121788 289836 251824 289864
rect 121788 289824 121794 289836
rect 251818 289824 251824 289836
rect 251876 289824 251882 289876
rect 121454 289756 121460 289808
rect 121512 289796 121518 289808
rect 124306 289796 124312 289808
rect 121512 289768 124312 289796
rect 121512 289756 121518 289768
rect 124306 289756 124312 289768
rect 124364 289756 124370 289808
rect 119798 289076 119804 289128
rect 119856 289116 119862 289128
rect 580258 289116 580264 289128
rect 119856 289088 580264 289116
rect 119856 289076 119862 289088
rect 580258 289076 580264 289088
rect 580316 289076 580322 289128
rect 121454 288328 121460 288380
rect 121512 288368 121518 288380
rect 133966 288368 133972 288380
rect 121512 288340 133972 288368
rect 121512 288328 121518 288340
rect 133966 288328 133972 288340
rect 134024 288368 134030 288380
rect 135162 288368 135168 288380
rect 134024 288340 135168 288368
rect 134024 288328 134030 288340
rect 135162 288328 135168 288340
rect 135220 288328 135226 288380
rect 135162 287648 135168 287700
rect 135220 287688 135226 287700
rect 582926 287688 582932 287700
rect 135220 287660 582932 287688
rect 135220 287648 135226 287660
rect 582926 287648 582932 287660
rect 582984 287648 582990 287700
rect 121730 287036 121736 287088
rect 121788 287076 121794 287088
rect 345014 287076 345020 287088
rect 121788 287048 345020 287076
rect 121788 287036 121794 287048
rect 345014 287036 345020 287048
rect 345072 287036 345078 287088
rect 65978 286968 65984 287020
rect 66036 287008 66042 287020
rect 67726 287008 67732 287020
rect 66036 286980 67732 287008
rect 66036 286968 66042 286980
rect 67726 286968 67732 286980
rect 67784 286968 67790 287020
rect 121454 286968 121460 287020
rect 121512 287008 121518 287020
rect 127066 287008 127072 287020
rect 121512 286980 127072 287008
rect 121512 286968 121518 286980
rect 127066 286968 127072 286980
rect 127124 286968 127130 287020
rect 120902 286356 120908 286408
rect 120960 286396 120966 286408
rect 136818 286396 136824 286408
rect 120960 286368 136824 286396
rect 120960 286356 120966 286368
rect 136818 286356 136824 286368
rect 136876 286356 136882 286408
rect 122282 286288 122288 286340
rect 122340 286328 122346 286340
rect 328730 286328 328736 286340
rect 122340 286300 328736 286328
rect 122340 286288 122346 286300
rect 328730 286288 328736 286300
rect 328788 286288 328794 286340
rect 120810 285676 120816 285728
rect 120868 285716 120874 285728
rect 177298 285716 177304 285728
rect 120868 285688 177304 285716
rect 120868 285676 120874 285688
rect 177298 285676 177304 285688
rect 177356 285676 177362 285728
rect 66070 285608 66076 285660
rect 66128 285648 66134 285660
rect 68186 285648 68192 285660
rect 66128 285620 68192 285648
rect 66128 285608 66134 285620
rect 68186 285608 68192 285620
rect 68244 285608 68250 285660
rect 121730 285608 121736 285660
rect 121788 285648 121794 285660
rect 125778 285648 125784 285660
rect 121788 285620 125784 285648
rect 121788 285608 121794 285620
rect 125778 285608 125784 285620
rect 125836 285608 125842 285660
rect 121546 284316 121552 284368
rect 121604 284356 121610 284368
rect 311158 284356 311164 284368
rect 121604 284328 311164 284356
rect 121604 284316 121610 284328
rect 311158 284316 311164 284328
rect 311216 284316 311222 284368
rect 60642 284248 60648 284300
rect 60700 284288 60706 284300
rect 67634 284288 67640 284300
rect 60700 284260 67640 284288
rect 60700 284248 60706 284260
rect 67634 284248 67640 284260
rect 67692 284248 67698 284300
rect 121454 284248 121460 284300
rect 121512 284288 121518 284300
rect 128538 284288 128544 284300
rect 121512 284260 128544 284288
rect 121512 284248 121518 284260
rect 128538 284248 128544 284260
rect 128596 284248 128602 284300
rect 121454 282888 121460 282940
rect 121512 282928 121518 282940
rect 325694 282928 325700 282940
rect 121512 282900 325700 282928
rect 121512 282888 121518 282900
rect 325694 282888 325700 282900
rect 325752 282888 325758 282940
rect 57790 282820 57796 282872
rect 57848 282860 57854 282872
rect 67634 282860 67640 282872
rect 57848 282832 67640 282860
rect 57848 282820 57854 282832
rect 67634 282820 67640 282832
rect 67692 282820 67698 282872
rect 121454 281528 121460 281580
rect 121512 281568 121518 281580
rect 240870 281568 240876 281580
rect 121512 281540 240876 281568
rect 121512 281528 121518 281540
rect 240870 281528 240876 281540
rect 240928 281528 240934 281580
rect 121454 280236 121460 280288
rect 121512 280276 121518 280288
rect 227070 280276 227076 280288
rect 121512 280248 227076 280276
rect 121512 280236 121518 280248
rect 227070 280236 227076 280248
rect 227128 280236 227134 280288
rect 52178 280168 52184 280220
rect 52236 280208 52242 280220
rect 67634 280208 67640 280220
rect 52236 280180 67640 280208
rect 52236 280168 52242 280180
rect 67634 280168 67640 280180
rect 67692 280168 67698 280220
rect 121546 280168 121552 280220
rect 121604 280208 121610 280220
rect 247770 280208 247776 280220
rect 121604 280180 247776 280208
rect 121604 280168 121610 280180
rect 247770 280168 247776 280180
rect 247828 280168 247834 280220
rect 46750 280100 46756 280152
rect 46808 280140 46814 280152
rect 67726 280140 67732 280152
rect 46808 280112 67732 280140
rect 46808 280100 46814 280112
rect 67726 280100 67732 280112
rect 67784 280100 67790 280152
rect 59262 280032 59268 280084
rect 59320 280072 59326 280084
rect 67634 280072 67640 280084
rect 59320 280044 67640 280072
rect 59320 280032 59326 280044
rect 67634 280032 67640 280044
rect 67692 280032 67698 280084
rect 25498 279420 25504 279472
rect 25556 279460 25562 279472
rect 46750 279460 46756 279472
rect 25556 279432 46756 279460
rect 25556 279420 25562 279432
rect 46750 279420 46756 279432
rect 46808 279420 46814 279472
rect 121730 279420 121736 279472
rect 121788 279460 121794 279472
rect 255314 279460 255320 279472
rect 121788 279432 255320 279460
rect 121788 279420 121794 279432
rect 255314 279420 255320 279432
rect 255372 279420 255378 279472
rect 121454 278808 121460 278860
rect 121512 278848 121518 278860
rect 148318 278848 148324 278860
rect 121512 278820 148324 278848
rect 121512 278808 121518 278820
rect 148318 278808 148324 278820
rect 148376 278808 148382 278860
rect 121546 278740 121552 278792
rect 121604 278780 121610 278792
rect 312538 278780 312544 278792
rect 121604 278752 312544 278780
rect 121604 278740 121610 278752
rect 312538 278740 312544 278752
rect 312596 278740 312602 278792
rect 48038 277448 48044 277500
rect 48096 277488 48102 277500
rect 67634 277488 67640 277500
rect 48096 277460 67640 277488
rect 48096 277448 48102 277460
rect 67634 277448 67640 277460
rect 67692 277448 67698 277500
rect 121454 277448 121460 277500
rect 121512 277488 121518 277500
rect 315298 277488 315304 277500
rect 121512 277460 315304 277488
rect 121512 277448 121518 277460
rect 315298 277448 315304 277460
rect 315356 277448 315362 277500
rect 46842 277380 46848 277432
rect 46900 277420 46906 277432
rect 67726 277420 67732 277432
rect 46900 277392 67732 277420
rect 46900 277380 46906 277392
rect 67726 277380 67732 277392
rect 67784 277380 67790 277432
rect 121546 277380 121552 277432
rect 121604 277420 121610 277432
rect 322198 277420 322204 277432
rect 121604 277392 322204 277420
rect 121604 277380 121610 277392
rect 322198 277380 322204 277392
rect 322256 277380 322262 277432
rect 121454 277312 121460 277364
rect 121512 277352 121518 277364
rect 129918 277352 129924 277364
rect 121512 277324 129924 277352
rect 121512 277312 121518 277324
rect 129918 277312 129924 277324
rect 129976 277312 129982 277364
rect 129918 276632 129924 276684
rect 129976 276672 129982 276684
rect 144086 276672 144092 276684
rect 129976 276644 144092 276672
rect 129976 276632 129982 276644
rect 144086 276632 144092 276644
rect 144144 276632 144150 276684
rect 50798 276088 50804 276140
rect 50856 276128 50862 276140
rect 67634 276128 67640 276140
rect 50856 276100 67640 276128
rect 50856 276088 50862 276100
rect 67634 276088 67640 276100
rect 67692 276088 67698 276140
rect 121454 276020 121460 276072
rect 121512 276060 121518 276072
rect 338206 276060 338212 276072
rect 121512 276032 338212 276060
rect 121512 276020 121518 276032
rect 338206 276020 338212 276032
rect 338264 276020 338270 276072
rect 64598 274728 64604 274780
rect 64656 274768 64662 274780
rect 67634 274768 67640 274780
rect 64656 274740 67640 274768
rect 64656 274728 64662 274740
rect 67634 274728 67640 274740
rect 67692 274728 67698 274780
rect 57790 274660 57796 274712
rect 57848 274700 57854 274712
rect 67818 274700 67824 274712
rect 57848 274672 67824 274700
rect 57848 274660 57854 274672
rect 67818 274660 67824 274672
rect 67876 274660 67882 274712
rect 44082 274592 44088 274644
rect 44140 274632 44146 274644
rect 67726 274632 67732 274644
rect 44140 274604 67732 274632
rect 44140 274592 44146 274604
rect 67726 274592 67732 274604
rect 67784 274592 67790 274644
rect 121454 274592 121460 274644
rect 121512 274632 121518 274644
rect 124858 274632 124864 274644
rect 121512 274604 124864 274632
rect 121512 274592 121518 274604
rect 124858 274592 124864 274604
rect 124916 274592 124922 274644
rect 121638 273912 121644 273964
rect 121696 273952 121702 273964
rect 468478 273952 468484 273964
rect 121696 273924 468484 273952
rect 121696 273912 121702 273924
rect 468478 273912 468484 273924
rect 468536 273912 468542 273964
rect 121454 273232 121460 273284
rect 121512 273272 121518 273284
rect 214558 273272 214564 273284
rect 121512 273244 214564 273272
rect 121512 273232 121518 273244
rect 214558 273232 214564 273244
rect 214616 273232 214622 273284
rect 121546 273164 121552 273216
rect 121604 273204 121610 273216
rect 125870 273204 125876 273216
rect 121604 273176 125876 273204
rect 121604 273164 121610 273176
rect 125870 273164 125876 273176
rect 125928 273164 125934 273216
rect 139394 273164 139400 273216
rect 139452 273204 139458 273216
rect 580166 273204 580172 273216
rect 139452 273176 580172 273204
rect 139452 273164 139458 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 124950 272484 124956 272536
rect 125008 272524 125014 272536
rect 139394 272524 139400 272536
rect 125008 272496 139400 272524
rect 125008 272484 125014 272496
rect 139394 272484 139400 272496
rect 139452 272484 139458 272536
rect 60274 271940 60280 271992
rect 60332 271980 60338 271992
rect 67634 271980 67640 271992
rect 60332 271952 67640 271980
rect 60332 271940 60338 271952
rect 67634 271940 67640 271952
rect 67692 271940 67698 271992
rect 59262 271872 59268 271924
rect 59320 271912 59326 271924
rect 67818 271912 67824 271924
rect 59320 271884 67824 271912
rect 59320 271872 59326 271884
rect 67818 271872 67824 271884
rect 67876 271872 67882 271924
rect 60550 271804 60556 271856
rect 60608 271844 60614 271856
rect 67726 271844 67732 271856
rect 60608 271816 67732 271844
rect 60608 271804 60614 271816
rect 67726 271804 67732 271816
rect 67784 271804 67790 271856
rect 61746 270512 61752 270564
rect 61804 270552 61810 270564
rect 67634 270552 67640 270564
rect 61804 270524 67640 270552
rect 61804 270512 61810 270524
rect 67634 270512 67640 270524
rect 67692 270512 67698 270564
rect 121454 270512 121460 270564
rect 121512 270552 121518 270564
rect 252646 270552 252652 270564
rect 121512 270524 252652 270552
rect 121512 270512 121518 270524
rect 252646 270512 252652 270524
rect 252704 270512 252710 270564
rect 144086 269764 144092 269816
rect 144144 269804 144150 269816
rect 580534 269804 580540 269816
rect 144144 269776 580540 269804
rect 144144 269764 144150 269776
rect 580534 269764 580540 269776
rect 580592 269764 580598 269816
rect 54754 269152 54760 269204
rect 54812 269192 54818 269204
rect 67726 269192 67732 269204
rect 54812 269164 67732 269192
rect 54812 269152 54818 269164
rect 67726 269152 67732 269164
rect 67784 269152 67790 269204
rect 53650 269084 53656 269136
rect 53708 269124 53714 269136
rect 67634 269124 67640 269136
rect 53708 269096 67640 269124
rect 53708 269084 53714 269096
rect 67634 269084 67640 269096
rect 67692 269084 67698 269136
rect 121454 269084 121460 269136
rect 121512 269124 121518 269136
rect 233878 269124 233884 269136
rect 121512 269096 233884 269124
rect 121512 269084 121518 269096
rect 233878 269084 233884 269096
rect 233936 269084 233942 269136
rect 121546 269016 121552 269068
rect 121604 269056 121610 269068
rect 132586 269056 132592 269068
rect 121604 269028 132592 269056
rect 121604 269016 121610 269028
rect 132586 269016 132592 269028
rect 132644 269016 132650 269068
rect 43990 268336 43996 268388
rect 44048 268376 44054 268388
rect 67634 268376 67640 268388
rect 44048 268348 67640 268376
rect 44048 268336 44054 268348
rect 67634 268336 67640 268348
rect 67692 268336 67698 268388
rect 121638 268336 121644 268388
rect 121696 268376 121702 268388
rect 252554 268376 252560 268388
rect 121696 268348 252560 268376
rect 121696 268336 121702 268348
rect 252554 268336 252560 268348
rect 252612 268336 252618 268388
rect 66162 268200 66168 268252
rect 66220 268240 66226 268252
rect 68186 268240 68192 268252
rect 66220 268212 68192 268240
rect 66220 268200 66226 268212
rect 68186 268200 68192 268212
rect 68244 268200 68250 268252
rect 43438 268064 43444 268116
rect 43496 268104 43502 268116
rect 43990 268104 43996 268116
rect 43496 268076 43996 268104
rect 43496 268064 43502 268076
rect 43990 268064 43996 268076
rect 44048 268064 44054 268116
rect 121454 267724 121460 267776
rect 121512 267764 121518 267776
rect 339494 267764 339500 267776
rect 121512 267736 339500 267764
rect 121512 267724 121518 267736
rect 339494 267724 339500 267736
rect 339552 267724 339558 267776
rect 41322 267656 41328 267708
rect 41380 267696 41386 267708
rect 67726 267696 67732 267708
rect 41380 267668 67732 267696
rect 41380 267656 41386 267668
rect 67726 267656 67732 267668
rect 67784 267656 67790 267708
rect 54938 267588 54944 267640
rect 54996 267628 55002 267640
rect 67634 267628 67640 267640
rect 54996 267600 67640 267628
rect 54996 267588 55002 267600
rect 67634 267588 67640 267600
rect 67692 267588 67698 267640
rect 3326 267112 3332 267164
rect 3384 267152 3390 267164
rect 7558 267152 7564 267164
rect 3384 267124 7564 267152
rect 3384 267112 3390 267124
rect 7558 267112 7564 267124
rect 7616 267112 7622 267164
rect 121454 266432 121460 266484
rect 121512 266472 121518 266484
rect 334066 266472 334072 266484
rect 121512 266444 334072 266472
rect 121512 266432 121518 266444
rect 334066 266432 334072 266444
rect 334124 266432 334130 266484
rect 121546 266364 121552 266416
rect 121604 266404 121610 266416
rect 347958 266404 347964 266416
rect 121604 266376 347964 266404
rect 121604 266364 121610 266376
rect 347958 266364 347964 266376
rect 348016 266364 348022 266416
rect 53558 266296 53564 266348
rect 53616 266336 53622 266348
rect 67634 266336 67640 266348
rect 53616 266308 67640 266336
rect 53616 266296 53622 266308
rect 67634 266296 67640 266308
rect 67692 266296 67698 266348
rect 125042 265616 125048 265668
rect 125100 265656 125106 265668
rect 580442 265656 580448 265668
rect 125100 265628 580448 265656
rect 125100 265616 125106 265628
rect 580442 265616 580448 265628
rect 580500 265616 580506 265668
rect 121454 265004 121460 265056
rect 121512 265044 121518 265056
rect 308490 265044 308496 265056
rect 121512 265016 308496 265044
rect 121512 265004 121518 265016
rect 308490 265004 308496 265016
rect 308548 265004 308554 265056
rect 56226 264936 56232 264988
rect 56284 264976 56290 264988
rect 67726 264976 67732 264988
rect 56284 264948 67732 264976
rect 56284 264936 56290 264948
rect 67726 264936 67732 264948
rect 67784 264936 67790 264988
rect 121546 264936 121552 264988
rect 121604 264976 121610 264988
rect 346486 264976 346492 264988
rect 121604 264948 346492 264976
rect 121604 264936 121610 264948
rect 346486 264936 346492 264948
rect 346544 264936 346550 264988
rect 48130 264868 48136 264920
rect 48188 264908 48194 264920
rect 67634 264908 67640 264920
rect 48188 264880 67640 264908
rect 48188 264868 48194 264880
rect 67634 264868 67640 264880
rect 67692 264868 67698 264920
rect 121454 264868 121460 264920
rect 121512 264908 121518 264920
rect 125686 264908 125692 264920
rect 121512 264880 125692 264908
rect 121512 264868 121518 264880
rect 125686 264868 125692 264880
rect 125744 264868 125750 264920
rect 18598 264188 18604 264240
rect 18656 264228 18662 264240
rect 48130 264228 48136 264240
rect 18656 264200 48136 264228
rect 18656 264188 18662 264200
rect 48130 264188 48136 264200
rect 48188 264188 48194 264240
rect 49510 263576 49516 263628
rect 49568 263616 49574 263628
rect 67726 263616 67732 263628
rect 49568 263588 67732 263616
rect 49568 263576 49574 263588
rect 67726 263576 67732 263588
rect 67784 263576 67790 263628
rect 121546 263576 121552 263628
rect 121604 263616 121610 263628
rect 233970 263616 233976 263628
rect 121604 263588 233976 263616
rect 121604 263576 121610 263588
rect 233970 263576 233976 263588
rect 234028 263576 234034 263628
rect 50890 263508 50896 263560
rect 50948 263548 50954 263560
rect 67634 263548 67640 263560
rect 50948 263520 67640 263548
rect 50948 263508 50954 263520
rect 67634 263508 67640 263520
rect 67692 263508 67698 263560
rect 121454 263508 121460 263560
rect 121512 263548 121518 263560
rect 123110 263548 123116 263560
rect 121512 263520 123116 263548
rect 121512 263508 121518 263520
rect 123110 263508 123116 263520
rect 123168 263508 123174 263560
rect 59078 262216 59084 262268
rect 59136 262256 59142 262268
rect 67634 262256 67640 262268
rect 59136 262228 67640 262256
rect 59136 262216 59142 262228
rect 67634 262216 67640 262228
rect 67692 262216 67698 262268
rect 121454 262216 121460 262268
rect 121512 262256 121518 262268
rect 338390 262256 338396 262268
rect 121512 262228 338396 262256
rect 121512 262216 121518 262228
rect 338390 262216 338396 262228
rect 338448 262216 338454 262268
rect 54846 260924 54852 260976
rect 54904 260964 54910 260976
rect 67634 260964 67640 260976
rect 54904 260936 67640 260964
rect 54904 260924 54910 260936
rect 67634 260924 67640 260936
rect 67692 260924 67698 260976
rect 53558 260856 53564 260908
rect 53616 260896 53622 260908
rect 67726 260896 67732 260908
rect 53616 260868 67732 260896
rect 53616 260856 53622 260868
rect 67726 260856 67732 260868
rect 67784 260856 67790 260908
rect 121546 260856 121552 260908
rect 121604 260896 121610 260908
rect 307110 260896 307116 260908
rect 121604 260868 307116 260896
rect 121604 260856 121610 260868
rect 307110 260856 307116 260868
rect 307168 260856 307174 260908
rect 61930 260788 61936 260840
rect 61988 260828 61994 260840
rect 67634 260828 67640 260840
rect 61988 260800 67640 260828
rect 61988 260788 61994 260800
rect 67634 260788 67640 260800
rect 67692 260788 67698 260840
rect 121454 260788 121460 260840
rect 121512 260828 121518 260840
rect 142154 260828 142160 260840
rect 121512 260800 142160 260828
rect 121512 260788 121518 260800
rect 142154 260788 142160 260800
rect 142212 260828 142218 260840
rect 143442 260828 143448 260840
rect 142212 260800 143448 260828
rect 142212 260788 142218 260800
rect 143442 260788 143448 260800
rect 143500 260788 143506 260840
rect 143442 260108 143448 260160
rect 143500 260148 143506 260160
rect 464338 260148 464344 260160
rect 143500 260120 464344 260148
rect 143500 260108 143506 260120
rect 464338 260108 464344 260120
rect 464396 260108 464402 260160
rect 61378 259428 61384 259480
rect 61436 259468 61442 259480
rect 67634 259468 67640 259480
rect 61436 259440 67640 259468
rect 61436 259428 61442 259440
rect 67634 259428 67640 259440
rect 67692 259428 67698 259480
rect 121454 259428 121460 259480
rect 121512 259468 121518 259480
rect 235258 259468 235264 259480
rect 121512 259440 235264 259468
rect 121512 259428 121518 259440
rect 235258 259428 235264 259440
rect 235316 259428 235322 259480
rect 121546 259360 121552 259412
rect 121604 259400 121610 259412
rect 132494 259400 132500 259412
rect 121604 259372 132500 259400
rect 121604 259360 121610 259372
rect 132494 259360 132500 259372
rect 132552 259360 132558 259412
rect 273898 259360 273904 259412
rect 273956 259400 273962 259412
rect 579890 259400 579896 259412
rect 273956 259372 579896 259400
rect 273956 259360 273962 259372
rect 579890 259360 579896 259372
rect 579948 259360 579954 259412
rect 60366 258136 60372 258188
rect 60424 258176 60430 258188
rect 67634 258176 67640 258188
rect 60424 258148 67640 258176
rect 60424 258136 60430 258148
rect 67634 258136 67640 258148
rect 67692 258136 67698 258188
rect 56410 258068 56416 258120
rect 56468 258108 56474 258120
rect 67726 258108 67732 258120
rect 56468 258080 67732 258108
rect 56468 258068 56474 258080
rect 67726 258068 67732 258080
rect 67784 258068 67790 258120
rect 121638 258068 121644 258120
rect 121696 258108 121702 258120
rect 347866 258108 347872 258120
rect 121696 258080 347872 258108
rect 121696 258068 121702 258080
rect 347866 258068 347872 258080
rect 347924 258068 347930 258120
rect 34330 258000 34336 258052
rect 34388 258040 34394 258052
rect 67634 258040 67640 258052
rect 34388 258012 67640 258040
rect 34388 258000 34394 258012
rect 67634 258000 67640 258012
rect 67692 258000 67698 258052
rect 121454 258000 121460 258052
rect 121512 258040 121518 258052
rect 128998 258040 129004 258052
rect 121512 258012 129004 258040
rect 121512 258000 121518 258012
rect 128998 258000 129004 258012
rect 129056 258000 129062 258052
rect 63310 257388 63316 257440
rect 63368 257428 63374 257440
rect 68370 257428 68376 257440
rect 63368 257400 68376 257428
rect 63368 257388 63374 257400
rect 68370 257388 68376 257400
rect 68428 257388 68434 257440
rect 4798 257320 4804 257372
rect 4856 257360 4862 257372
rect 34330 257360 34336 257372
rect 4856 257332 34336 257360
rect 4856 257320 4862 257332
rect 34330 257320 34336 257332
rect 34388 257320 34394 257372
rect 60642 257320 60648 257372
rect 60700 257360 60706 257372
rect 68278 257360 68284 257372
rect 60700 257332 68284 257360
rect 60700 257320 60706 257332
rect 68278 257320 68284 257332
rect 68336 257320 68342 257372
rect 63218 256708 63224 256760
rect 63276 256748 63282 256760
rect 67634 256748 67640 256760
rect 63276 256720 67640 256748
rect 63276 256708 63282 256720
rect 67634 256708 67640 256720
rect 67692 256708 67698 256760
rect 121546 256708 121552 256760
rect 121604 256748 121610 256760
rect 220078 256748 220084 256760
rect 121604 256720 220084 256748
rect 121604 256708 121610 256720
rect 220078 256708 220084 256720
rect 220136 256708 220142 256760
rect 121454 256640 121460 256692
rect 121512 256680 121518 256692
rect 129826 256680 129832 256692
rect 121512 256652 129832 256680
rect 121512 256640 121518 256652
rect 129826 256640 129832 256652
rect 129884 256640 129890 256692
rect 121546 256572 121552 256624
rect 121604 256612 121610 256624
rect 126974 256612 126980 256624
rect 121604 256584 126980 256612
rect 121604 256572 121610 256584
rect 126974 256572 126980 256584
rect 127032 256572 127038 256624
rect 120902 255960 120908 256012
rect 120960 256000 120966 256012
rect 580350 256000 580356 256012
rect 120960 255972 580356 256000
rect 120960 255960 120966 255972
rect 580350 255960 580356 255972
rect 580408 255960 580414 256012
rect 3142 255212 3148 255264
rect 3200 255252 3206 255264
rect 34882 255252 34888 255264
rect 3200 255224 34888 255252
rect 3200 255212 3206 255224
rect 34882 255212 34888 255224
rect 34940 255212 34946 255264
rect 55122 255212 55128 255264
rect 55180 255252 55186 255264
rect 67634 255252 67640 255264
rect 55180 255224 67640 255252
rect 55180 255212 55186 255224
rect 67634 255212 67640 255224
rect 67692 255212 67698 255264
rect 56318 254600 56324 254652
rect 56376 254640 56382 254652
rect 61654 254640 61660 254652
rect 56376 254612 61660 254640
rect 56376 254600 56382 254612
rect 61654 254600 61660 254612
rect 61712 254640 61718 254652
rect 67634 254640 67640 254652
rect 61712 254612 67640 254640
rect 61712 254600 61718 254612
rect 67634 254600 67640 254612
rect 67692 254600 67698 254652
rect 34882 254532 34888 254584
rect 34940 254572 34946 254584
rect 35802 254572 35808 254584
rect 34940 254544 35808 254572
rect 34940 254532 34946 254544
rect 35802 254532 35808 254544
rect 35860 254572 35866 254584
rect 58618 254572 58624 254584
rect 35860 254544 58624 254572
rect 35860 254532 35866 254544
rect 58618 254532 58624 254544
rect 58676 254532 58682 254584
rect 121454 253988 121460 254040
rect 121512 254028 121518 254040
rect 246390 254028 246396 254040
rect 121512 254000 246396 254028
rect 121512 253988 121518 254000
rect 246390 253988 246396 254000
rect 246448 253988 246454 254040
rect 121546 253920 121552 253972
rect 121604 253960 121610 253972
rect 314010 253960 314016 253972
rect 121604 253932 314016 253960
rect 121604 253920 121610 253932
rect 314010 253920 314016 253932
rect 314068 253920 314074 253972
rect 54478 253852 54484 253904
rect 54536 253892 54542 253904
rect 56502 253892 56508 253904
rect 54536 253864 56508 253892
rect 54536 253852 54542 253864
rect 56502 253852 56508 253864
rect 56560 253892 56566 253904
rect 67634 253892 67640 253904
rect 56560 253864 67640 253892
rect 56560 253852 56566 253864
rect 67634 253852 67640 253864
rect 67692 253852 67698 253904
rect 121546 252628 121552 252680
rect 121604 252668 121610 252680
rect 263594 252668 263600 252680
rect 121604 252640 263600 252668
rect 121604 252628 121610 252640
rect 263594 252628 263600 252640
rect 263652 252628 263658 252680
rect 64506 252560 64512 252612
rect 64564 252600 64570 252612
rect 67634 252600 67640 252612
rect 64564 252572 67640 252600
rect 64564 252560 64570 252572
rect 67634 252560 67640 252572
rect 67692 252560 67698 252612
rect 121454 252560 121460 252612
rect 121512 252600 121518 252612
rect 350718 252600 350724 252612
rect 121512 252572 350724 252600
rect 121512 252560 121518 252572
rect 350718 252560 350724 252572
rect 350776 252560 350782 252612
rect 64690 251268 64696 251320
rect 64748 251308 64754 251320
rect 67726 251308 67732 251320
rect 64748 251280 67732 251308
rect 64748 251268 64754 251280
rect 67726 251268 67732 251280
rect 67784 251268 67790 251320
rect 56502 251200 56508 251252
rect 56560 251240 56566 251252
rect 67634 251240 67640 251252
rect 56560 251212 67640 251240
rect 56560 251200 56566 251212
rect 67634 251200 67640 251212
rect 67692 251200 67698 251252
rect 121454 251200 121460 251252
rect 121512 251240 121518 251252
rect 331306 251240 331312 251252
rect 121512 251212 331312 251240
rect 121512 251200 121518 251212
rect 331306 251200 331312 251212
rect 331364 251200 331370 251252
rect 120442 250996 120448 251048
rect 120500 251036 120506 251048
rect 123018 251036 123024 251048
rect 120500 251008 123024 251036
rect 120500 250996 120506 251008
rect 123018 250996 123024 251008
rect 123076 250996 123082 251048
rect 65886 249840 65892 249892
rect 65944 249880 65950 249892
rect 67634 249880 67640 249892
rect 65944 249852 67640 249880
rect 65944 249840 65950 249852
rect 67634 249840 67640 249852
rect 67692 249840 67698 249892
rect 57606 249772 57612 249824
rect 57664 249812 57670 249824
rect 67726 249812 67732 249824
rect 57664 249784 67732 249812
rect 57664 249772 57670 249784
rect 67726 249772 67732 249784
rect 67784 249772 67790 249824
rect 121546 249772 121552 249824
rect 121604 249812 121610 249824
rect 238110 249812 238116 249824
rect 121604 249784 238116 249812
rect 121604 249772 121610 249784
rect 238110 249772 238116 249784
rect 238168 249772 238174 249824
rect 49602 249704 49608 249756
rect 49660 249744 49666 249756
rect 67634 249744 67640 249756
rect 49660 249716 67640 249744
rect 49660 249704 49666 249716
rect 67634 249704 67640 249716
rect 67692 249704 67698 249756
rect 121454 249704 121460 249756
rect 121512 249744 121518 249756
rect 140866 249744 140872 249756
rect 121512 249716 140872 249744
rect 121512 249704 121518 249716
rect 140866 249704 140872 249716
rect 140924 249704 140930 249756
rect 59170 249636 59176 249688
rect 59228 249676 59234 249688
rect 61378 249676 61384 249688
rect 59228 249648 61384 249676
rect 59228 249636 59234 249648
rect 61378 249636 61384 249648
rect 61436 249636 61442 249688
rect 120718 249500 120724 249552
rect 120776 249540 120782 249552
rect 121454 249540 121460 249552
rect 120776 249512 121460 249540
rect 120776 249500 120782 249512
rect 121454 249500 121460 249512
rect 121512 249500 121518 249552
rect 66070 248616 66076 248668
rect 66128 248656 66134 248668
rect 68094 248656 68100 248668
rect 66128 248628 68100 248656
rect 66128 248616 66134 248628
rect 68094 248616 68100 248628
rect 68152 248616 68158 248668
rect 121546 248412 121552 248464
rect 121604 248452 121610 248464
rect 210418 248452 210424 248464
rect 121604 248424 210424 248452
rect 121604 248412 121610 248424
rect 210418 248412 210424 248424
rect 210476 248412 210482 248464
rect 121454 248344 121460 248396
rect 121512 248344 121518 248396
rect 121638 248344 121644 248396
rect 121696 248384 121702 248396
rect 147674 248384 147680 248396
rect 121696 248356 147680 248384
rect 121696 248344 121702 248356
rect 147674 248344 147680 248356
rect 147732 248344 147738 248396
rect 121472 248316 121500 248344
rect 121730 248316 121736 248328
rect 121472 248288 121736 248316
rect 121730 248276 121736 248288
rect 121788 248276 121794 248328
rect 177298 247664 177304 247716
rect 177356 247704 177362 247716
rect 580350 247704 580356 247716
rect 177356 247676 580356 247704
rect 177356 247664 177362 247676
rect 580350 247664 580356 247676
rect 580408 247664 580414 247716
rect 62022 247120 62028 247172
rect 62080 247160 62086 247172
rect 67726 247160 67732 247172
rect 62080 247132 67732 247160
rect 62080 247120 62086 247132
rect 67726 247120 67732 247132
rect 67784 247120 67790 247172
rect 61930 247052 61936 247104
rect 61988 247092 61994 247104
rect 67634 247092 67640 247104
rect 61988 247064 67640 247092
rect 61988 247052 61994 247064
rect 67634 247052 67640 247064
rect 67692 247052 67698 247104
rect 121454 247052 121460 247104
rect 121512 247092 121518 247104
rect 266354 247092 266360 247104
rect 121512 247064 266360 247092
rect 121512 247052 121518 247064
rect 266354 247052 266360 247064
rect 266412 247052 266418 247104
rect 121546 245692 121552 245744
rect 121604 245732 121610 245744
rect 224310 245732 224316 245744
rect 121604 245704 224316 245732
rect 121604 245692 121610 245704
rect 224310 245692 224316 245704
rect 224368 245692 224374 245744
rect 121454 245624 121460 245676
rect 121512 245664 121518 245676
rect 231210 245664 231216 245676
rect 121512 245636 231216 245664
rect 121512 245624 121518 245636
rect 231210 245624 231216 245636
rect 231268 245624 231274 245676
rect 61838 245556 61844 245608
rect 61896 245596 61902 245608
rect 67634 245596 67640 245608
rect 61896 245568 67640 245596
rect 61896 245556 61902 245568
rect 67634 245556 67640 245568
rect 67692 245556 67698 245608
rect 65978 244264 65984 244316
rect 66036 244304 66042 244316
rect 68094 244304 68100 244316
rect 66036 244276 68100 244304
rect 66036 244264 66042 244276
rect 68094 244264 68100 244276
rect 68152 244264 68158 244316
rect 342438 244264 342444 244316
rect 342496 244304 342502 244316
rect 580166 244304 580172 244316
rect 342496 244276 580172 244304
rect 342496 244264 342502 244276
rect 580166 244264 580172 244276
rect 580224 244264 580230 244316
rect 11698 244196 11704 244248
rect 11756 244236 11762 244248
rect 39850 244236 39856 244248
rect 11756 244208 39856 244236
rect 11756 244196 11762 244208
rect 39850 244196 39856 244208
rect 39908 244236 39914 244248
rect 67634 244236 67640 244248
rect 39908 244208 67640 244236
rect 39908 244196 39914 244208
rect 67634 244196 67640 244208
rect 67692 244196 67698 244248
rect 121454 244196 121460 244248
rect 121512 244236 121518 244248
rect 134058 244236 134064 244248
rect 121512 244208 134064 244236
rect 121512 244196 121518 244208
rect 134058 244196 134064 244208
rect 134116 244196 134122 244248
rect 121638 243516 121644 243568
rect 121696 243556 121702 243568
rect 321554 243556 321560 243568
rect 121696 243528 321560 243556
rect 121696 243516 121702 243528
rect 321554 243516 321560 243528
rect 321612 243516 321618 243568
rect 121546 242904 121552 242956
rect 121604 242944 121610 242956
rect 335538 242944 335544 242956
rect 121604 242916 335544 242944
rect 121604 242904 121610 242916
rect 335538 242904 335544 242916
rect 335596 242904 335602 242956
rect 121454 242836 121460 242888
rect 121512 242876 121518 242888
rect 132678 242876 132684 242888
rect 121512 242848 132684 242876
rect 121512 242836 121518 242848
rect 132678 242836 132684 242848
rect 132736 242876 132742 242888
rect 342438 242876 342444 242888
rect 132736 242848 342444 242876
rect 132736 242836 132742 242848
rect 342438 242836 342444 242848
rect 342496 242836 342502 242888
rect 121546 242768 121552 242820
rect 121604 242808 121610 242820
rect 128446 242808 128452 242820
rect 121604 242780 128452 242808
rect 121604 242768 121610 242780
rect 128446 242768 128452 242780
rect 128504 242768 128510 242820
rect 63402 241476 63408 241528
rect 63460 241516 63466 241528
rect 67634 241516 67640 241528
rect 63460 241488 67640 241516
rect 63460 241476 63466 241488
rect 67634 241476 67640 241488
rect 67692 241476 67698 241528
rect 121454 241476 121460 241528
rect 121512 241516 121518 241528
rect 249794 241516 249800 241528
rect 121512 241488 249800 241516
rect 121512 241476 121518 241488
rect 249794 241476 249800 241488
rect 249852 241476 249858 241528
rect 121546 240728 121552 240780
rect 121604 240768 121610 240780
rect 135254 240768 135260 240780
rect 121604 240740 135260 240768
rect 121604 240728 121610 240740
rect 135254 240728 135260 240740
rect 135312 240728 135318 240780
rect 3050 240116 3056 240168
rect 3108 240156 3114 240168
rect 11146 240156 11152 240168
rect 3108 240128 11152 240156
rect 3108 240116 3114 240128
rect 11146 240116 11152 240128
rect 11204 240116 11210 240168
rect 119890 240116 119896 240168
rect 119948 240156 119954 240168
rect 329834 240156 329840 240168
rect 119948 240128 329840 240156
rect 119948 240116 119954 240128
rect 329834 240116 329840 240128
rect 329892 240116 329898 240168
rect 65886 239912 65892 239964
rect 65944 239952 65950 239964
rect 72510 239952 72516 239964
rect 65944 239924 72516 239952
rect 65944 239912 65950 239924
rect 72510 239912 72516 239924
rect 72568 239912 72574 239964
rect 75914 239776 75920 239828
rect 75972 239816 75978 239828
rect 77098 239816 77104 239828
rect 75972 239788 77104 239816
rect 75972 239776 75978 239788
rect 77098 239776 77104 239788
rect 77156 239776 77162 239828
rect 78674 239776 78680 239828
rect 78732 239816 78738 239828
rect 79674 239816 79680 239828
rect 78732 239788 79680 239816
rect 78732 239776 78738 239788
rect 79674 239776 79680 239788
rect 79732 239776 79738 239828
rect 86954 239776 86960 239828
rect 87012 239816 87018 239828
rect 88046 239816 88052 239828
rect 87012 239788 88052 239816
rect 87012 239776 87018 239788
rect 88046 239776 88052 239788
rect 88104 239776 88110 239828
rect 89714 239776 89720 239828
rect 89772 239816 89778 239828
rect 90622 239816 90628 239828
rect 89772 239788 90628 239816
rect 89772 239776 89778 239788
rect 90622 239776 90628 239788
rect 90680 239776 90686 239828
rect 100754 239776 100760 239828
rect 100812 239816 100818 239828
rect 101570 239816 101576 239828
rect 100812 239788 101576 239816
rect 100812 239776 100818 239788
rect 101570 239776 101576 239788
rect 101628 239776 101634 239828
rect 103606 239776 103612 239828
rect 103664 239816 103670 239828
rect 104790 239816 104796 239828
rect 103664 239788 104796 239816
rect 103664 239776 103670 239788
rect 104790 239776 104796 239788
rect 104848 239776 104854 239828
rect 104894 239776 104900 239828
rect 104952 239816 104958 239828
rect 106078 239816 106084 239828
rect 104952 239788 106084 239816
rect 104952 239776 104958 239788
rect 106078 239776 106084 239788
rect 106136 239776 106142 239828
rect 107654 239776 107660 239828
rect 107712 239816 107718 239828
rect 108654 239816 108660 239828
rect 107712 239788 108660 239816
rect 107712 239776 107718 239788
rect 108654 239776 108660 239788
rect 108712 239776 108718 239828
rect 114554 239776 114560 239828
rect 114612 239816 114618 239828
rect 115738 239816 115744 239828
rect 114612 239788 115744 239816
rect 114612 239776 114618 239788
rect 115738 239776 115744 239788
rect 115796 239776 115802 239828
rect 121454 239708 121460 239760
rect 121512 239748 121518 239760
rect 124858 239748 124864 239760
rect 121512 239720 124864 239748
rect 121512 239708 121518 239720
rect 124858 239708 124864 239720
rect 124916 239708 124922 239760
rect 69750 239504 69756 239556
rect 69808 239544 69814 239556
rect 83550 239544 83556 239556
rect 69808 239516 83556 239544
rect 69808 239504 69814 239516
rect 83550 239504 83556 239516
rect 83608 239504 83614 239556
rect 64506 239436 64512 239488
rect 64564 239476 64570 239488
rect 339586 239476 339592 239488
rect 64564 239448 339592 239476
rect 64564 239436 64570 239448
rect 339586 239436 339592 239448
rect 339644 239436 339650 239488
rect 63218 239368 63224 239420
rect 63276 239408 63282 239420
rect 342438 239408 342444 239420
rect 63276 239380 342444 239408
rect 63276 239368 63282 239380
rect 342438 239368 342444 239380
rect 342496 239368 342502 239420
rect 84286 239300 84292 239352
rect 84344 239340 84350 239352
rect 85482 239340 85488 239352
rect 84344 239312 85488 239340
rect 84344 239300 84350 239312
rect 85482 239300 85488 239312
rect 85540 239300 85546 239352
rect 99006 238960 99012 239012
rect 99064 239000 99070 239012
rect 131114 239000 131120 239012
rect 99064 238972 131120 239000
rect 99064 238960 99070 238972
rect 131114 238960 131120 238972
rect 131172 238960 131178 239012
rect 115106 238892 115112 238944
rect 115164 238932 115170 238944
rect 124214 238932 124220 238944
rect 115164 238904 124220 238932
rect 115164 238892 115170 238904
rect 124214 238892 124220 238904
rect 124272 238892 124278 238944
rect 114462 238824 114468 238876
rect 114520 238864 114526 238876
rect 127158 238864 127164 238876
rect 114520 238836 127164 238864
rect 114520 238824 114526 238836
rect 127158 238824 127164 238836
rect 127216 238824 127222 238876
rect 52362 238756 52368 238808
rect 52420 238796 52426 238808
rect 95786 238796 95792 238808
rect 52420 238768 95792 238796
rect 52420 238756 52426 238768
rect 95786 238756 95792 238768
rect 95844 238756 95850 238808
rect 7558 238688 7564 238740
rect 7616 238728 7622 238740
rect 57698 238728 57704 238740
rect 7616 238700 57704 238728
rect 7616 238688 7622 238700
rect 57698 238688 57704 238700
rect 57756 238728 57762 238740
rect 86770 238728 86776 238740
rect 57756 238700 86776 238728
rect 57756 238688 57762 238700
rect 86770 238688 86776 238700
rect 86828 238688 86834 238740
rect 89346 238688 89352 238740
rect 89404 238728 89410 238740
rect 129734 238728 129740 238740
rect 89404 238700 129740 238728
rect 89404 238688 89410 238700
rect 129734 238688 129740 238700
rect 129792 238688 129798 238740
rect 48222 238620 48228 238672
rect 48280 238660 48286 238672
rect 82262 238660 82268 238672
rect 48280 238632 82268 238660
rect 48280 238620 48286 238632
rect 82262 238620 82268 238632
rect 82320 238620 82326 238672
rect 91922 238620 91928 238672
rect 91980 238660 91986 238672
rect 120902 238660 120908 238672
rect 91980 238632 120908 238660
rect 91980 238620 91986 238632
rect 120902 238620 120908 238632
rect 120960 238620 120966 238672
rect 63126 238552 63132 238604
rect 63184 238592 63190 238604
rect 72602 238592 72608 238604
rect 63184 238564 72608 238592
rect 63184 238552 63190 238564
rect 72602 238552 72608 238564
rect 72660 238552 72666 238604
rect 118326 238552 118332 238604
rect 118384 238592 118390 238604
rect 136726 238592 136732 238604
rect 118384 238564 136732 238592
rect 118384 238552 118390 238564
rect 136726 238552 136732 238564
rect 136784 238552 136790 238604
rect 106734 238484 106740 238536
rect 106792 238524 106798 238536
rect 121454 238524 121460 238536
rect 106792 238496 121460 238524
rect 106792 238484 106798 238496
rect 121454 238484 121460 238496
rect 121512 238484 121518 238536
rect 102870 238144 102876 238196
rect 102928 238184 102934 238196
rect 106918 238184 106924 238196
rect 102928 238156 106924 238184
rect 102928 238144 102934 238156
rect 106918 238144 106924 238156
rect 106976 238144 106982 238196
rect 82906 238076 82912 238128
rect 82964 238116 82970 238128
rect 88978 238116 88984 238128
rect 82964 238088 88984 238116
rect 82964 238076 82970 238088
rect 88978 238076 88984 238088
rect 89036 238076 89042 238128
rect 96430 238076 96436 238128
rect 96488 238116 96494 238128
rect 184198 238116 184204 238128
rect 96488 238088 184204 238116
rect 96488 238076 96494 238088
rect 184198 238076 184204 238088
rect 184256 238076 184262 238128
rect 68830 238008 68836 238060
rect 68888 238048 68894 238060
rect 327166 238048 327172 238060
rect 68888 238020 327172 238048
rect 68888 238008 68894 238020
rect 327166 238008 327172 238020
rect 327224 238008 327230 238060
rect 71314 237464 71320 237516
rect 71372 237504 71378 237516
rect 75178 237504 75184 237516
rect 71372 237476 75184 237504
rect 71372 237464 71378 237476
rect 75178 237464 75184 237476
rect 75236 237464 75242 237516
rect 69934 237396 69940 237448
rect 69992 237436 69998 237448
rect 72418 237436 72424 237448
rect 69992 237408 72424 237436
rect 69992 237396 69998 237408
rect 72418 237396 72424 237408
rect 72476 237396 72482 237448
rect 75822 237328 75828 237380
rect 75880 237368 75886 237380
rect 143534 237368 143540 237380
rect 75880 237340 143540 237368
rect 75880 237328 75886 237340
rect 143534 237328 143540 237340
rect 143592 237328 143598 237380
rect 68922 236648 68928 236700
rect 68980 236688 68986 236700
rect 286318 236688 286324 236700
rect 68980 236660 286324 236688
rect 68980 236648 68986 236660
rect 286318 236648 286324 236660
rect 286376 236648 286382 236700
rect 324958 236648 324964 236700
rect 325016 236688 325022 236700
rect 347774 236688 347780 236700
rect 325016 236660 347780 236688
rect 325016 236648 325022 236660
rect 347774 236648 347780 236660
rect 347832 236648 347838 236700
rect 11146 235900 11152 235952
rect 11204 235940 11210 235952
rect 37090 235940 37096 235952
rect 11204 235912 37096 235940
rect 11204 235900 11210 235912
rect 37090 235900 37096 235912
rect 37148 235940 37154 235952
rect 103514 235940 103520 235952
rect 37148 235912 103520 235940
rect 37148 235900 37154 235912
rect 103514 235900 103520 235912
rect 103572 235900 103578 235952
rect 117682 235900 117688 235952
rect 117740 235940 117746 235952
rect 133874 235940 133880 235952
rect 117740 235912 133880 235940
rect 117740 235900 117746 235912
rect 133874 235900 133880 235912
rect 133932 235940 133938 235952
rect 135162 235940 135168 235952
rect 133932 235912 135168 235940
rect 133932 235900 133938 235912
rect 135162 235900 135168 235912
rect 135220 235900 135226 235952
rect 58618 235832 58624 235884
rect 58676 235872 58682 235884
rect 112530 235872 112536 235884
rect 58676 235844 112536 235872
rect 58676 235832 58682 235844
rect 112530 235832 112536 235844
rect 112588 235832 112594 235884
rect 53742 235764 53748 235816
rect 53800 235804 53806 235816
rect 107378 235804 107384 235816
rect 53800 235776 107384 235804
rect 53800 235764 53806 235776
rect 107378 235764 107384 235776
rect 107436 235764 107442 235816
rect 52270 235696 52276 235748
rect 52328 235736 52334 235748
rect 76558 235736 76564 235748
rect 52328 235708 76564 235736
rect 52328 235696 52334 235708
rect 76558 235696 76564 235708
rect 76616 235696 76622 235748
rect 81618 235696 81624 235748
rect 81676 235736 81682 235748
rect 120810 235736 120816 235748
rect 81676 235708 120816 235736
rect 81676 235696 81682 235708
rect 120810 235696 120816 235708
rect 120868 235696 120874 235748
rect 91278 235628 91284 235680
rect 91336 235668 91342 235680
rect 124950 235668 124956 235680
rect 91336 235640 124956 235668
rect 91336 235628 91342 235640
rect 124950 235628 124956 235640
rect 125008 235628 125014 235680
rect 135162 235220 135168 235272
rect 135220 235260 135226 235272
rect 180150 235260 180156 235272
rect 135220 235232 180156 235260
rect 135220 235220 135226 235232
rect 180150 235220 180156 235232
rect 180208 235220 180214 235272
rect 45462 234540 45468 234592
rect 45520 234580 45526 234592
rect 109034 234580 109040 234592
rect 45520 234552 109040 234580
rect 45520 234540 45526 234552
rect 109034 234540 109040 234552
rect 109092 234540 109098 234592
rect 110598 234540 110604 234592
rect 110656 234580 110662 234592
rect 111058 234580 111064 234592
rect 110656 234552 111064 234580
rect 110656 234540 110662 234552
rect 111058 234540 111064 234552
rect 111116 234580 111122 234592
rect 136634 234580 136640 234592
rect 111116 234552 136640 234580
rect 111116 234540 111122 234552
rect 136634 234540 136640 234552
rect 136692 234540 136698 234592
rect 88978 234472 88984 234524
rect 89036 234512 89042 234524
rect 128354 234512 128360 234524
rect 89036 234484 128360 234512
rect 89036 234472 89042 234484
rect 128354 234472 128360 234484
rect 128412 234472 128418 234524
rect 109034 234132 109040 234184
rect 109092 234172 109098 234184
rect 109954 234172 109960 234184
rect 109092 234144 109960 234172
rect 109092 234132 109098 234144
rect 109954 234132 109960 234144
rect 110012 234132 110018 234184
rect 80330 233928 80336 233980
rect 80388 233968 80394 233980
rect 320910 233968 320916 233980
rect 80388 233940 320916 233968
rect 80388 233928 80394 233940
rect 320910 233928 320916 233940
rect 320968 233928 320974 233980
rect 128354 233860 128360 233912
rect 128412 233900 128418 233912
rect 582742 233900 582748 233912
rect 128412 233872 582748 233900
rect 128412 233860 128418 233872
rect 582742 233860 582748 233872
rect 582800 233860 582806 233912
rect 84102 231820 84108 231872
rect 84160 231860 84166 231872
rect 84838 231860 84844 231872
rect 84160 231832 84844 231860
rect 84160 231820 84166 231832
rect 84838 231820 84844 231832
rect 84896 231820 84902 231872
rect 64598 231140 64604 231192
rect 64656 231180 64662 231192
rect 133138 231180 133144 231192
rect 64656 231152 133144 231180
rect 64656 231140 64662 231152
rect 133138 231140 133144 231152
rect 133196 231140 133202 231192
rect 78306 231072 78312 231124
rect 78364 231112 78370 231124
rect 267734 231112 267740 231124
rect 78364 231084 267740 231112
rect 78364 231072 78370 231084
rect 267734 231072 267740 231084
rect 267792 231072 267798 231124
rect 60182 230392 60188 230444
rect 60240 230432 60246 230444
rect 60458 230432 60464 230444
rect 60240 230404 60464 230432
rect 60240 230392 60246 230404
rect 60458 230392 60464 230404
rect 60516 230432 60522 230444
rect 83366 230432 83372 230444
rect 60516 230404 83372 230432
rect 60516 230392 60522 230404
rect 83366 230392 83372 230404
rect 83424 230392 83430 230444
rect 17218 229712 17224 229764
rect 17276 229752 17282 229764
rect 60182 229752 60188 229764
rect 17276 229724 60188 229752
rect 17276 229712 17282 229724
rect 60182 229712 60188 229724
rect 60240 229712 60246 229764
rect 72510 229712 72516 229764
rect 72568 229752 72574 229764
rect 336734 229752 336740 229764
rect 72568 229724 336740 229752
rect 72568 229712 72574 229724
rect 336734 229712 336740 229724
rect 336792 229712 336798 229764
rect 97626 228420 97632 228472
rect 97684 228460 97690 228472
rect 333974 228460 333980 228472
rect 97684 228432 333980 228460
rect 97684 228420 97690 228432
rect 333974 228420 333980 228432
rect 334032 228420 334038 228472
rect 88334 228352 88340 228404
rect 88392 228392 88398 228404
rect 353386 228392 353392 228404
rect 88392 228364 353392 228392
rect 88392 228352 88398 228364
rect 353386 228352 353392 228364
rect 353444 228352 353450 228404
rect 63402 226992 63408 227044
rect 63460 227032 63466 227044
rect 214650 227032 214656 227044
rect 63460 227004 214656 227032
rect 63460 226992 63466 227004
rect 214650 226992 214656 227004
rect 214708 226992 214714 227044
rect 3602 225564 3608 225616
rect 3660 225604 3666 225616
rect 120074 225604 120080 225616
rect 3660 225576 120080 225604
rect 3660 225564 3666 225576
rect 120074 225564 120080 225576
rect 120132 225564 120138 225616
rect 78766 224272 78772 224324
rect 78824 224312 78830 224324
rect 228358 224312 228364 224324
rect 78824 224284 228364 224312
rect 78824 224272 78830 224284
rect 228358 224272 228364 224284
rect 228416 224272 228422 224324
rect 95050 224204 95056 224256
rect 95108 224244 95114 224256
rect 345106 224244 345112 224256
rect 95108 224216 345112 224244
rect 95108 224204 95114 224216
rect 345106 224204 345112 224216
rect 345164 224204 345170 224256
rect 75178 221484 75184 221536
rect 75236 221524 75242 221536
rect 242158 221524 242164 221536
rect 75236 221496 242164 221524
rect 75236 221484 75242 221496
rect 242158 221484 242164 221496
rect 242216 221484 242222 221536
rect 56226 221416 56232 221468
rect 56284 221456 56290 221468
rect 340874 221456 340880 221468
rect 56284 221428 340880 221456
rect 56284 221416 56290 221428
rect 340874 221416 340880 221428
rect 340932 221416 340938 221468
rect 114554 220124 114560 220176
rect 114612 220164 114618 220176
rect 311250 220164 311256 220176
rect 114612 220136 311256 220164
rect 114612 220124 114618 220136
rect 311250 220124 311256 220136
rect 311308 220124 311314 220176
rect 46842 220056 46848 220108
rect 46900 220096 46906 220108
rect 296070 220096 296076 220108
rect 46900 220068 296076 220096
rect 46900 220056 46906 220068
rect 296070 220056 296076 220068
rect 296128 220056 296134 220108
rect 110414 218764 110420 218816
rect 110472 218804 110478 218816
rect 256970 218804 256976 218816
rect 110472 218776 256976 218804
rect 110472 218764 110478 218776
rect 256970 218764 256976 218776
rect 257028 218764 257034 218816
rect 103606 218696 103612 218748
rect 103664 218736 103670 218748
rect 325786 218736 325792 218748
rect 103664 218708 325792 218736
rect 103664 218696 103670 218708
rect 325786 218696 325792 218708
rect 325844 218696 325850 218748
rect 82078 217268 82084 217320
rect 82136 217308 82142 217320
rect 300210 217308 300216 217320
rect 82136 217280 300216 217308
rect 82136 217268 82142 217280
rect 300210 217268 300216 217280
rect 300268 217268 300274 217320
rect 99466 215976 99472 216028
rect 99524 216016 99530 216028
rect 253934 216016 253940 216028
rect 99524 215988 253940 216016
rect 99524 215976 99530 215988
rect 253934 215976 253940 215988
rect 253992 215976 253998 216028
rect 93946 215908 93952 215960
rect 94004 215948 94010 215960
rect 322934 215948 322940 215960
rect 94004 215920 322940 215948
rect 94004 215908 94010 215920
rect 322934 215908 322940 215920
rect 322992 215908 322998 215960
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 18598 215268 18604 215280
rect 3384 215240 18604 215268
rect 3384 215228 3390 215240
rect 18598 215228 18604 215240
rect 18656 215228 18662 215280
rect 56410 214616 56416 214668
rect 56468 214656 56474 214668
rect 280154 214656 280160 214668
rect 56468 214628 280160 214656
rect 56468 214616 56474 214628
rect 280154 214616 280160 214628
rect 280212 214616 280218 214668
rect 103698 214548 103704 214600
rect 103756 214588 103762 214600
rect 352098 214588 352104 214600
rect 103756 214560 352104 214588
rect 103756 214548 103762 214560
rect 352098 214548 352104 214560
rect 352156 214548 352162 214600
rect 89806 213324 89812 213376
rect 89864 213364 89870 213376
rect 254118 213364 254124 213376
rect 89864 213336 254124 213364
rect 89864 213324 89870 213336
rect 254118 213324 254124 213336
rect 254176 213324 254182 213376
rect 87046 213256 87052 213308
rect 87104 213296 87110 213308
rect 327074 213296 327080 213308
rect 87104 213268 327080 213296
rect 87104 213256 87110 213268
rect 327074 213256 327080 213268
rect 327132 213256 327138 213308
rect 54846 213188 54852 213240
rect 54904 213228 54910 213240
rect 316678 213228 316684 213240
rect 54904 213200 316684 213228
rect 54904 213188 54910 213200
rect 316678 213188 316684 213200
rect 316736 213188 316742 213240
rect 104986 211760 104992 211812
rect 105044 211800 105050 211812
rect 331490 211800 331496 211812
rect 105044 211772 331496 211800
rect 105044 211760 105050 211772
rect 331490 211760 331496 211772
rect 331548 211760 331554 211812
rect 61930 210468 61936 210520
rect 61988 210508 61994 210520
rect 236638 210508 236644 210520
rect 61988 210480 236644 210508
rect 61988 210468 61994 210480
rect 236638 210468 236644 210480
rect 236696 210468 236702 210520
rect 83458 210400 83464 210452
rect 83516 210440 83522 210452
rect 335446 210440 335452 210452
rect 83516 210412 335452 210440
rect 83516 210400 83522 210412
rect 335446 210400 335452 210412
rect 335504 210400 335510 210452
rect 100846 209176 100852 209228
rect 100904 209216 100910 209228
rect 254026 209216 254032 209228
rect 100904 209188 254032 209216
rect 100904 209176 100910 209188
rect 254026 209176 254032 209188
rect 254084 209176 254090 209228
rect 48038 209108 48044 209160
rect 48096 209148 48102 209160
rect 270494 209148 270500 209160
rect 48096 209120 270500 209148
rect 48096 209108 48102 209120
rect 270494 209108 270500 209120
rect 270552 209108 270558 209160
rect 113174 209040 113180 209092
rect 113232 209080 113238 209092
rect 338298 209080 338304 209092
rect 113232 209052 338304 209080
rect 113232 209040 113238 209052
rect 338298 209040 338304 209052
rect 338356 209040 338362 209092
rect 86954 207680 86960 207732
rect 87012 207720 87018 207732
rect 252830 207720 252836 207732
rect 87012 207692 252836 207720
rect 87012 207680 87018 207692
rect 252830 207680 252836 207692
rect 252888 207680 252894 207732
rect 74626 207612 74632 207664
rect 74684 207652 74690 207664
rect 278866 207652 278872 207664
rect 74684 207624 278872 207652
rect 74684 207612 74690 207624
rect 278866 207612 278872 207624
rect 278924 207612 278930 207664
rect 111794 206252 111800 206304
rect 111852 206292 111858 206304
rect 255406 206292 255412 206304
rect 111852 206264 255412 206292
rect 111852 206252 111858 206264
rect 255406 206252 255412 206264
rect 255464 206252 255470 206304
rect 89714 204960 89720 205012
rect 89772 205000 89778 205012
rect 281626 205000 281632 205012
rect 89772 204972 281632 205000
rect 89772 204960 89778 204972
rect 281626 204960 281632 204972
rect 281684 204960 281690 205012
rect 59078 204892 59084 204944
rect 59136 204932 59142 204944
rect 259454 204932 259460 204944
rect 59136 204904 259460 204932
rect 59136 204892 59142 204904
rect 259454 204892 259460 204904
rect 259512 204892 259518 204944
rect 50798 203532 50804 203584
rect 50856 203572 50862 203584
rect 263778 203572 263784 203584
rect 50856 203544 263784 203572
rect 50856 203532 50862 203544
rect 263778 203532 263784 203544
rect 263836 203532 263842 203584
rect 106918 202240 106924 202292
rect 106976 202280 106982 202292
rect 239398 202280 239404 202292
rect 106976 202252 239404 202280
rect 106976 202240 106982 202252
rect 239398 202240 239404 202252
rect 239456 202240 239462 202292
rect 100754 202172 100760 202224
rect 100812 202212 100818 202224
rect 252738 202212 252744 202224
rect 100812 202184 252744 202212
rect 100812 202172 100818 202184
rect 252738 202172 252744 202184
rect 252796 202172 252802 202224
rect 72418 202104 72424 202156
rect 72476 202144 72482 202156
rect 343910 202144 343916 202156
rect 72476 202116 343916 202144
rect 72476 202104 72482 202116
rect 343910 202104 343916 202116
rect 343968 202104 343974 202156
rect 93854 200880 93860 200932
rect 93912 200920 93918 200932
rect 255498 200920 255504 200932
rect 93912 200892 255504 200920
rect 93912 200880 93918 200892
rect 255498 200880 255504 200892
rect 255556 200880 255562 200932
rect 96614 200812 96620 200864
rect 96672 200852 96678 200864
rect 260834 200852 260840 200864
rect 96672 200824 260840 200852
rect 96672 200812 96678 200824
rect 260834 200812 260840 200824
rect 260892 200812 260898 200864
rect 107746 200744 107752 200796
rect 107804 200784 107810 200796
rect 328638 200784 328644 200796
rect 107804 200756 328644 200784
rect 107804 200744 107810 200756
rect 328638 200744 328644 200756
rect 328696 200744 328702 200796
rect 133138 199520 133144 199572
rect 133196 199560 133202 199572
rect 265066 199560 265072 199572
rect 133196 199532 265072 199560
rect 133196 199520 133202 199532
rect 265066 199520 265072 199532
rect 265124 199520 265130 199572
rect 115934 199452 115940 199504
rect 115992 199492 115998 199504
rect 270678 199492 270684 199504
rect 115992 199464 270684 199492
rect 115992 199452 115998 199464
rect 270678 199452 270684 199464
rect 270736 199452 270742 199504
rect 77294 199384 77300 199436
rect 77352 199424 77358 199436
rect 329926 199424 329932 199436
rect 77352 199396 329932 199424
rect 77352 199384 77358 199396
rect 329926 199384 329932 199396
rect 329984 199384 329990 199436
rect 251818 198160 251824 198212
rect 251876 198200 251882 198212
rect 274818 198200 274824 198212
rect 251876 198172 274824 198200
rect 251876 198160 251882 198172
rect 274818 198160 274824 198172
rect 274876 198160 274882 198212
rect 60274 198092 60280 198144
rect 60332 198132 60338 198144
rect 272058 198132 272064 198144
rect 60332 198104 272064 198132
rect 60332 198092 60338 198104
rect 272058 198092 272064 198104
rect 272116 198092 272122 198144
rect 92566 198024 92572 198076
rect 92624 198064 92630 198076
rect 330018 198064 330024 198076
rect 92624 198036 330024 198064
rect 92624 198024 92630 198036
rect 330018 198024 330024 198036
rect 330076 198024 330082 198076
rect 76558 197956 76564 198008
rect 76616 197996 76622 198008
rect 582834 197996 582840 198008
rect 76616 197968 582840 197996
rect 76616 197956 76622 197968
rect 582834 197956 582840 197968
rect 582892 197956 582898 198008
rect 92474 196732 92480 196784
rect 92532 196772 92538 196784
rect 261018 196772 261024 196784
rect 92532 196744 261024 196772
rect 92532 196732 92538 196744
rect 261018 196732 261024 196744
rect 261076 196732 261082 196784
rect 69014 196664 69020 196716
rect 69072 196704 69078 196716
rect 251174 196704 251180 196716
rect 69072 196676 251180 196704
rect 69072 196664 69078 196676
rect 251174 196664 251180 196676
rect 251232 196664 251238 196716
rect 107654 196596 107660 196648
rect 107712 196636 107718 196648
rect 328546 196636 328552 196648
rect 107712 196608 328552 196636
rect 107712 196596 107718 196608
rect 328546 196596 328552 196608
rect 328604 196596 328610 196648
rect 54754 195372 54760 195424
rect 54812 195412 54818 195424
rect 269206 195412 269212 195424
rect 54812 195384 269212 195412
rect 54812 195372 54818 195384
rect 269206 195372 269212 195384
rect 269264 195372 269270 195424
rect 124858 195304 124864 195356
rect 124916 195344 124922 195356
rect 345198 195344 345204 195356
rect 124916 195316 345204 195344
rect 124916 195304 124922 195316
rect 345198 195304 345204 195316
rect 345256 195304 345262 195356
rect 86218 195236 86224 195288
rect 86276 195276 86282 195288
rect 582650 195276 582656 195288
rect 86276 195248 582656 195276
rect 86276 195236 86282 195248
rect 582650 195236 582656 195248
rect 582708 195236 582714 195288
rect 247770 194012 247776 194064
rect 247828 194052 247834 194064
rect 340966 194052 340972 194064
rect 247828 194024 340972 194052
rect 247828 194012 247834 194024
rect 340966 194012 340972 194024
rect 341024 194012 341030 194064
rect 142798 193944 142804 193996
rect 142856 193984 142862 193996
rect 259730 193984 259736 193996
rect 142856 193956 259736 193984
rect 142856 193944 142862 193956
rect 259730 193944 259736 193956
rect 259788 193944 259794 193996
rect 57606 193876 57612 193928
rect 57664 193916 57670 193928
rect 273346 193916 273352 193928
rect 57664 193888 273352 193916
rect 57664 193876 57670 193888
rect 273346 193876 273352 193888
rect 273404 193876 273410 193928
rect 78674 193808 78680 193860
rect 78732 193848 78738 193860
rect 335630 193848 335636 193860
rect 78732 193820 335636 193848
rect 78732 193808 78738 193820
rect 335630 193808 335636 193820
rect 335688 193808 335694 193860
rect 152458 192720 152464 192772
rect 152516 192760 152522 192772
rect 200758 192760 200764 192772
rect 152516 192732 200764 192760
rect 152516 192720 152522 192732
rect 200758 192720 200764 192732
rect 200816 192720 200822 192772
rect 146938 192652 146944 192704
rect 146996 192692 147002 192704
rect 209130 192692 209136 192704
rect 146996 192664 209136 192692
rect 146996 192652 147002 192664
rect 209130 192652 209136 192664
rect 209188 192652 209194 192704
rect 199378 192584 199384 192636
rect 199436 192624 199442 192636
rect 280246 192624 280252 192636
rect 199436 192596 280252 192624
rect 199436 192584 199442 192596
rect 280246 192584 280252 192596
rect 280304 192584 280310 192636
rect 84286 192516 84292 192568
rect 84344 192556 84350 192568
rect 254210 192556 254216 192568
rect 84344 192528 254216 192556
rect 84344 192516 84350 192528
rect 254210 192516 254216 192528
rect 254268 192516 254274 192568
rect 70394 192448 70400 192500
rect 70452 192488 70458 192500
rect 321738 192488 321744 192500
rect 70452 192460 321744 192488
rect 70452 192448 70458 192460
rect 321738 192448 321744 192460
rect 321796 192448 321802 192500
rect 148318 191292 148324 191344
rect 148376 191332 148382 191344
rect 239490 191332 239496 191344
rect 148376 191304 239496 191332
rect 148376 191292 148382 191304
rect 239490 191292 239496 191304
rect 239548 191292 239554 191344
rect 246298 191292 246304 191344
rect 246356 191332 246362 191344
rect 277486 191332 277492 191344
rect 246356 191304 277492 191332
rect 246356 191292 246362 191304
rect 277486 191292 277492 191304
rect 277544 191292 277550 191344
rect 192478 191224 192484 191276
rect 192536 191264 192542 191276
rect 331398 191264 331404 191276
rect 192536 191236 331404 191264
rect 192536 191224 192542 191236
rect 331398 191224 331404 191236
rect 331456 191224 331462 191276
rect 59262 191156 59268 191208
rect 59320 191196 59326 191208
rect 256786 191196 256792 191208
rect 59320 191168 256792 191196
rect 59320 191156 59326 191168
rect 256786 191156 256792 191168
rect 256844 191156 256850 191208
rect 62022 191088 62028 191140
rect 62080 191128 62086 191140
rect 262306 191128 262312 191140
rect 62080 191100 262312 191128
rect 62080 191088 62086 191100
rect 262306 191088 262312 191100
rect 262364 191088 262370 191140
rect 213270 189864 213276 189916
rect 213328 189904 213334 189916
rect 281718 189904 281724 189916
rect 213328 189876 281724 189904
rect 213328 189864 213334 189876
rect 281718 189864 281724 189876
rect 281776 189864 281782 189916
rect 144178 189796 144184 189848
rect 144236 189836 144242 189848
rect 242250 189836 242256 189848
rect 144236 189808 242256 189836
rect 144236 189796 144242 189808
rect 242250 189796 242256 189808
rect 242308 189796 242314 189848
rect 56502 189728 56508 189780
rect 56560 189768 56566 189780
rect 199470 189768 199476 189780
rect 56560 189740 199476 189768
rect 56560 189728 56566 189740
rect 199470 189728 199476 189740
rect 199528 189728 199534 189780
rect 249150 189728 249156 189780
rect 249208 189768 249214 189780
rect 336826 189768 336832 189780
rect 249208 189740 336832 189768
rect 249208 189728 249214 189740
rect 336826 189728 336832 189740
rect 336884 189728 336890 189780
rect 107562 189048 107568 189100
rect 107620 189088 107626 189100
rect 188430 189088 188436 189100
rect 107620 189060 188436 189088
rect 107620 189048 107626 189060
rect 188430 189048 188436 189060
rect 188488 189048 188494 189100
rect 209222 188640 209228 188692
rect 209280 188680 209286 188692
rect 261110 188680 261116 188692
rect 209280 188652 261116 188680
rect 209280 188640 209286 188652
rect 261110 188640 261116 188652
rect 261168 188640 261174 188692
rect 202230 188572 202236 188624
rect 202288 188612 202294 188624
rect 267918 188612 267924 188624
rect 202288 188584 267924 188612
rect 202288 188572 202294 188584
rect 267918 188572 267924 188584
rect 267976 188572 267982 188624
rect 15838 188504 15844 188556
rect 15896 188544 15902 188556
rect 109034 188544 109040 188556
rect 15896 188516 109040 188544
rect 15896 188504 15902 188516
rect 109034 188504 109040 188516
rect 109092 188504 109098 188556
rect 141418 188504 141424 188556
rect 141476 188544 141482 188556
rect 262398 188544 262404 188556
rect 141476 188516 262404 188544
rect 141476 188504 141482 188516
rect 262398 188504 262404 188516
rect 262456 188504 262462 188556
rect 69198 188436 69204 188488
rect 69256 188476 69262 188488
rect 319622 188476 319628 188488
rect 69256 188448 319628 188476
rect 69256 188436 69262 188448
rect 319622 188436 319628 188448
rect 319680 188436 319686 188488
rect 69106 188368 69112 188420
rect 69164 188408 69170 188420
rect 341150 188408 341156 188420
rect 69164 188380 341156 188408
rect 69164 188368 69170 188380
rect 341150 188368 341156 188380
rect 341208 188368 341214 188420
rect 57790 188300 57796 188352
rect 57848 188340 57854 188352
rect 334250 188340 334256 188352
rect 57848 188312 334256 188340
rect 57848 188300 57854 188312
rect 334250 188300 334256 188312
rect 334308 188300 334314 188352
rect 129642 187756 129648 187808
rect 129700 187796 129706 187808
rect 177298 187796 177304 187808
rect 129700 187768 177304 187796
rect 129700 187756 129706 187768
rect 177298 187756 177304 187768
rect 177356 187756 177362 187808
rect 104802 187688 104808 187740
rect 104860 187728 104866 187740
rect 173250 187728 173256 187740
rect 104860 187700 173256 187728
rect 104860 187688 104866 187700
rect 173250 187688 173256 187700
rect 173308 187688 173314 187740
rect 203518 187008 203524 187060
rect 203576 187048 203582 187060
rect 276198 187048 276204 187060
rect 203576 187020 276204 187048
rect 203576 187008 203582 187020
rect 276198 187008 276204 187020
rect 276256 187008 276262 187060
rect 73246 186940 73252 186992
rect 73304 186980 73310 186992
rect 323118 186980 323124 186992
rect 73304 186952 323124 186980
rect 73304 186940 73310 186952
rect 323118 186940 323124 186952
rect 323176 186940 323182 186992
rect 100662 186464 100668 186516
rect 100720 186504 100726 186516
rect 169110 186504 169116 186516
rect 100720 186476 169116 186504
rect 100720 186464 100726 186476
rect 169110 186464 169116 186476
rect 169168 186464 169174 186516
rect 99282 186396 99288 186448
rect 99340 186436 99346 186448
rect 171778 186436 171784 186448
rect 99340 186408 171784 186436
rect 99340 186396 99346 186408
rect 171778 186396 171784 186408
rect 171836 186396 171842 186448
rect 119982 186328 119988 186380
rect 120040 186368 120046 186380
rect 214742 186368 214748 186380
rect 120040 186340 214748 186368
rect 120040 186328 120046 186340
rect 214742 186328 214748 186340
rect 214800 186328 214806 186380
rect 151078 185920 151084 185972
rect 151136 185960 151142 185972
rect 187050 185960 187056 185972
rect 151136 185932 187056 185960
rect 151136 185920 151142 185932
rect 187050 185920 187056 185932
rect 187108 185920 187114 185972
rect 232590 185920 232596 185972
rect 232648 185960 232654 185972
rect 266446 185960 266452 185972
rect 232648 185932 266452 185960
rect 232648 185920 232654 185932
rect 266446 185920 266452 185932
rect 266504 185920 266510 185972
rect 65978 185852 65984 185904
rect 66036 185892 66042 185904
rect 274726 185892 274732 185904
rect 66036 185864 274732 185892
rect 66036 185852 66042 185864
rect 274726 185852 274732 185864
rect 274784 185852 274790 185904
rect 99374 185784 99380 185836
rect 99432 185824 99438 185836
rect 325970 185824 325976 185836
rect 99432 185796 325976 185824
rect 99432 185784 99438 185796
rect 325970 185784 325976 185796
rect 326028 185784 326034 185836
rect 104894 185716 104900 185768
rect 104952 185756 104958 185768
rect 339678 185756 339684 185768
rect 104952 185728 339684 185756
rect 104952 185716 104958 185728
rect 339678 185716 339684 185728
rect 339736 185716 339742 185768
rect 80054 185648 80060 185700
rect 80112 185688 80118 185700
rect 327350 185688 327356 185700
rect 80112 185660 327356 185688
rect 80112 185648 80118 185660
rect 327350 185648 327356 185660
rect 327408 185648 327414 185700
rect 67450 185580 67456 185632
rect 67508 185620 67514 185632
rect 324314 185620 324320 185632
rect 67508 185592 324320 185620
rect 67508 185580 67514 185592
rect 324314 185580 324320 185592
rect 324372 185580 324378 185632
rect 214650 184356 214656 184408
rect 214708 184396 214714 184408
rect 270586 184396 270592 184408
rect 214708 184368 270592 184396
rect 214708 184356 214714 184368
rect 270586 184356 270592 184368
rect 270644 184356 270650 184408
rect 67542 184288 67548 184340
rect 67600 184328 67606 184340
rect 251266 184328 251272 184340
rect 67600 184300 251272 184328
rect 67600 184288 67606 184300
rect 251266 184288 251272 184300
rect 251324 184288 251330 184340
rect 73154 184220 73160 184272
rect 73212 184260 73218 184272
rect 323210 184260 323216 184272
rect 73212 184232 323216 184260
rect 73212 184220 73218 184232
rect 323210 184220 323216 184232
rect 323268 184220 323274 184272
rect 64690 184152 64696 184204
rect 64748 184192 64754 184204
rect 341058 184192 341064 184204
rect 64748 184164 341064 184192
rect 64748 184152 64754 184164
rect 341058 184152 341064 184164
rect 341116 184152 341122 184204
rect 128262 183608 128268 183660
rect 128320 183648 128326 183660
rect 166534 183648 166540 183660
rect 128320 183620 166540 183648
rect 128320 183608 128326 183620
rect 166534 183608 166540 183620
rect 166592 183608 166598 183660
rect 114462 183540 114468 183592
rect 114520 183580 114526 183592
rect 169294 183580 169300 183592
rect 114520 183552 169300 183580
rect 114520 183540 114526 183552
rect 169294 183540 169300 183552
rect 169352 183540 169358 183592
rect 224218 183132 224224 183184
rect 224276 183172 224282 183184
rect 258258 183172 258264 183184
rect 224276 183144 258264 183172
rect 224276 183132 224282 183144
rect 258258 183132 258264 183144
rect 258316 183132 258322 183184
rect 226978 183064 226984 183116
rect 227036 183104 227042 183116
rect 263870 183104 263876 183116
rect 227036 183076 263876 183104
rect 227036 183064 227042 183076
rect 263870 183064 263876 183076
rect 263928 183064 263934 183116
rect 155218 182996 155224 183048
rect 155276 183036 155282 183048
rect 193858 183036 193864 183048
rect 155276 183008 193864 183036
rect 155276 182996 155282 183008
rect 193858 182996 193864 183008
rect 193916 182996 193922 183048
rect 222838 182996 222844 183048
rect 222896 183036 222902 183048
rect 266538 183036 266544 183048
rect 222896 183008 266544 183036
rect 222896 182996 222902 183008
rect 266538 182996 266544 183008
rect 266596 182996 266602 183048
rect 311158 182996 311164 183048
rect 311216 183036 311222 183048
rect 332778 183036 332784 183048
rect 311216 183008 332784 183036
rect 311216 182996 311222 183008
rect 332778 182996 332784 183008
rect 332836 182996 332842 183048
rect 63310 182928 63316 182980
rect 63368 182968 63374 182980
rect 271966 182968 271972 182980
rect 63368 182940 271972 182968
rect 63368 182928 63374 182940
rect 271966 182928 271972 182940
rect 272024 182928 272030 182980
rect 307110 182928 307116 182980
rect 307168 182968 307174 182980
rect 334158 182968 334164 182980
rect 307168 182940 334164 182968
rect 307168 182928 307174 182940
rect 334158 182928 334164 182940
rect 334216 182928 334222 182980
rect 84194 182860 84200 182912
rect 84252 182900 84258 182912
rect 325878 182900 325884 182912
rect 84252 182872 325884 182900
rect 84252 182860 84258 182872
rect 325878 182860 325884 182872
rect 325936 182860 325942 182912
rect 75914 182792 75920 182844
rect 75972 182832 75978 182844
rect 321646 182832 321652 182844
rect 75972 182804 321652 182832
rect 75972 182792 75978 182804
rect 321646 182792 321652 182804
rect 321704 182792 321710 182844
rect 116946 182248 116952 182300
rect 117004 182288 117010 182300
rect 170582 182288 170588 182300
rect 117004 182260 170588 182288
rect 117004 182248 117010 182260
rect 170582 182248 170588 182260
rect 170640 182248 170646 182300
rect 110690 182180 110696 182232
rect 110748 182220 110754 182232
rect 167638 182220 167644 182232
rect 110748 182192 167644 182220
rect 110748 182180 110754 182192
rect 167638 182180 167644 182192
rect 167696 182180 167702 182232
rect 231210 181704 231216 181756
rect 231268 181744 231274 181756
rect 258074 181744 258080 181756
rect 231268 181716 258080 181744
rect 231268 181704 231274 181716
rect 258074 181704 258080 181716
rect 258132 181704 258138 181756
rect 238018 181636 238024 181688
rect 238076 181676 238082 181688
rect 264974 181676 264980 181688
rect 238076 181648 264980 181676
rect 238076 181636 238082 181648
rect 264974 181636 264980 181648
rect 265032 181636 265038 181688
rect 122098 181568 122104 181620
rect 122156 181608 122162 181620
rect 171134 181608 171140 181620
rect 122156 181580 171140 181608
rect 122156 181568 122162 181580
rect 171134 181568 171140 181580
rect 171192 181568 171198 181620
rect 207658 181568 207664 181620
rect 207716 181608 207722 181620
rect 273530 181608 273536 181620
rect 207716 181580 273536 181608
rect 207716 181568 207722 181580
rect 273530 181568 273536 181580
rect 273588 181568 273594 181620
rect 59170 181500 59176 181552
rect 59228 181540 59234 181552
rect 336918 181540 336924 181552
rect 59228 181512 336924 181540
rect 59228 181500 59234 181512
rect 336918 181500 336924 181512
rect 336976 181500 336982 181552
rect 53558 181432 53564 181484
rect 53616 181472 53622 181484
rect 345290 181472 345296 181484
rect 53616 181444 345296 181472
rect 53616 181432 53622 181444
rect 345290 181432 345296 181444
rect 345348 181432 345354 181484
rect 120902 180956 120908 181008
rect 120960 180996 120966 181008
rect 167730 180996 167736 181008
rect 120960 180968 167736 180996
rect 120960 180956 120966 180968
rect 167730 180956 167736 180968
rect 167788 180956 167794 181008
rect 115842 180888 115848 180940
rect 115900 180928 115906 180940
rect 166442 180928 166448 180940
rect 115900 180900 166448 180928
rect 115900 180888 115906 180900
rect 166442 180888 166448 180900
rect 166500 180888 166506 180940
rect 130746 180820 130752 180872
rect 130804 180860 130810 180872
rect 214650 180860 214656 180872
rect 130804 180832 214656 180860
rect 130804 180820 130810 180832
rect 214650 180820 214656 180832
rect 214708 180820 214714 180872
rect 239398 180412 239404 180464
rect 239456 180452 239462 180464
rect 258350 180452 258356 180464
rect 239456 180424 258356 180452
rect 239456 180412 239462 180424
rect 258350 180412 258356 180424
rect 258408 180412 258414 180464
rect 233970 180344 233976 180396
rect 234028 180384 234034 180396
rect 265250 180384 265256 180396
rect 234028 180356 265256 180384
rect 234028 180344 234034 180356
rect 265250 180344 265256 180356
rect 265308 180344 265314 180396
rect 166258 180276 166264 180328
rect 166316 180316 166322 180328
rect 182818 180316 182824 180328
rect 166316 180288 182824 180316
rect 166316 180276 166322 180288
rect 182818 180276 182824 180288
rect 182876 180276 182882 180328
rect 222930 180276 222936 180328
rect 222988 180316 222994 180328
rect 263686 180316 263692 180328
rect 222988 180288 263692 180316
rect 222988 180276 222994 180288
rect 263686 180276 263692 180288
rect 263744 180276 263750 180328
rect 160738 180208 160744 180260
rect 160796 180248 160802 180260
rect 192478 180248 192484 180260
rect 160796 180220 192484 180248
rect 160796 180208 160802 180220
rect 192478 180208 192484 180220
rect 192536 180208 192542 180260
rect 220078 180208 220084 180260
rect 220136 180248 220142 180260
rect 267826 180248 267832 180260
rect 220136 180220 267832 180248
rect 220136 180208 220142 180220
rect 267826 180208 267832 180220
rect 267884 180208 267890 180260
rect 66070 180140 66076 180192
rect 66128 180180 66134 180192
rect 273438 180180 273444 180192
rect 66128 180152 273444 180180
rect 66128 180140 66134 180152
rect 273438 180140 273444 180152
rect 273496 180140 273502 180192
rect 300118 180140 300124 180192
rect 300176 180180 300182 180192
rect 332594 180180 332600 180192
rect 300176 180152 332600 180180
rect 300176 180140 300182 180152
rect 332594 180140 332600 180152
rect 332652 180140 332658 180192
rect 71866 180072 71872 180124
rect 71924 180112 71930 180124
rect 327258 180112 327264 180124
rect 71924 180084 327264 180112
rect 71924 180072 71930 180084
rect 327258 180072 327264 180084
rect 327316 180072 327322 180124
rect 125410 179460 125416 179512
rect 125468 179500 125474 179512
rect 167914 179500 167920 179512
rect 125468 179472 167920 179500
rect 125468 179460 125474 179472
rect 167914 179460 167920 179472
rect 167972 179460 167978 179512
rect 112162 179392 112168 179444
rect 112220 179432 112226 179444
rect 170490 179432 170496 179444
rect 112220 179404 170496 179432
rect 112220 179392 112226 179404
rect 170490 179392 170496 179404
rect 170548 179392 170554 179444
rect 235258 178916 235264 178968
rect 235316 178956 235322 178968
rect 265158 178956 265164 178968
rect 235316 178928 265164 178956
rect 235316 178916 235322 178928
rect 265158 178916 265164 178928
rect 265216 178916 265222 178968
rect 227070 178848 227076 178900
rect 227128 178888 227134 178900
rect 259546 178888 259552 178900
rect 227128 178860 259552 178888
rect 227128 178848 227134 178860
rect 259546 178848 259552 178860
rect 259604 178848 259610 178900
rect 214558 178780 214564 178832
rect 214616 178820 214622 178832
rect 249334 178820 249340 178832
rect 214616 178792 249340 178820
rect 214616 178780 214622 178792
rect 249334 178780 249340 178792
rect 249392 178780 249398 178832
rect 315298 178780 315304 178832
rect 315356 178820 315362 178832
rect 339770 178820 339776 178832
rect 315356 178792 339776 178820
rect 315356 178780 315362 178792
rect 339770 178780 339776 178792
rect 339828 178780 339834 178832
rect 66162 178712 66168 178764
rect 66220 178752 66226 178764
rect 251358 178752 251364 178764
rect 66220 178724 251364 178752
rect 66220 178712 66226 178724
rect 251358 178712 251364 178724
rect 251416 178712 251422 178764
rect 311250 178712 311256 178764
rect 311308 178752 311314 178764
rect 342530 178752 342536 178764
rect 311308 178724 342536 178752
rect 311308 178712 311314 178724
rect 342530 178712 342536 178724
rect 342588 178712 342594 178764
rect 102134 178644 102140 178696
rect 102192 178684 102198 178696
rect 346578 178684 346584 178696
rect 102192 178656 346584 178684
rect 102192 178644 102198 178656
rect 346578 178644 346584 178656
rect 346636 178644 346642 178696
rect 133138 178236 133144 178288
rect 133196 178276 133202 178288
rect 164878 178276 164884 178288
rect 133196 178248 164884 178276
rect 133196 178236 133202 178248
rect 164878 178236 164884 178248
rect 164936 178236 164942 178288
rect 148226 178168 148232 178220
rect 148284 178208 148290 178220
rect 181438 178208 181444 178220
rect 148284 178180 181444 178208
rect 148284 178168 148290 178180
rect 181438 178168 181444 178180
rect 181496 178168 181502 178220
rect 123294 178100 123300 178152
rect 123352 178140 123358 178152
rect 166350 178140 166356 178152
rect 123352 178112 166356 178140
rect 123352 178100 123358 178112
rect 166350 178100 166356 178112
rect 166408 178100 166414 178152
rect 110046 178032 110052 178084
rect 110104 178072 110110 178084
rect 170398 178072 170404 178084
rect 110104 178044 170404 178072
rect 110104 178032 110110 178044
rect 170398 178032 170404 178044
rect 170456 178032 170462 178084
rect 272610 178032 272616 178084
rect 272668 178072 272674 178084
rect 316034 178072 316040 178084
rect 272668 178044 316040 178072
rect 272668 178032 272674 178044
rect 316034 178032 316040 178044
rect 316092 178032 316098 178084
rect 242158 177964 242164 178016
rect 242216 178004 242222 178016
rect 249886 178004 249892 178016
rect 242216 177976 249892 178004
rect 242216 177964 242222 177976
rect 249886 177964 249892 177976
rect 249944 177964 249950 178016
rect 247678 177556 247684 177608
rect 247736 177596 247742 177608
rect 258166 177596 258172 177608
rect 247736 177568 258172 177596
rect 247736 177556 247742 177568
rect 258166 177556 258172 177568
rect 258224 177556 258230 177608
rect 319530 177556 319536 177608
rect 319588 177596 319594 177608
rect 330110 177596 330116 177608
rect 319588 177568 330116 177596
rect 319588 177556 319594 177568
rect 330110 177556 330116 177568
rect 330168 177556 330174 177608
rect 233878 177488 233884 177540
rect 233936 177528 233942 177540
rect 260926 177528 260932 177540
rect 233936 177500 260932 177528
rect 233936 177488 233942 177500
rect 260926 177488 260932 177500
rect 260984 177488 260990 177540
rect 319622 177488 319628 177540
rect 319680 177528 319686 177540
rect 331214 177528 331220 177540
rect 319680 177500 331220 177528
rect 319680 177488 319686 177500
rect 331214 177488 331220 177500
rect 331272 177488 331278 177540
rect 228358 177420 228364 177472
rect 228416 177460 228422 177472
rect 259638 177460 259644 177472
rect 228416 177432 259644 177460
rect 228416 177420 228422 177432
rect 259638 177420 259644 177432
rect 259696 177420 259702 177472
rect 314010 177420 314016 177472
rect 314068 177460 314074 177472
rect 332686 177460 332692 177472
rect 314068 177432 332692 177460
rect 314068 177420 314074 177432
rect 332686 177420 332692 177432
rect 332744 177420 332750 177472
rect 224310 177352 224316 177404
rect 224368 177392 224374 177404
rect 262490 177392 262496 177404
rect 224368 177364 262496 177392
rect 224368 177352 224374 177364
rect 262490 177352 262496 177364
rect 262548 177352 262554 177404
rect 307018 177352 307024 177404
rect 307076 177392 307082 177404
rect 350534 177392 350540 177404
rect 307076 177364 350540 177392
rect 307076 177352 307082 177364
rect 350534 177352 350540 177364
rect 350592 177352 350598 177404
rect 184198 177284 184204 177336
rect 184256 177324 184262 177336
rect 324406 177324 324412 177336
rect 184256 177296 324412 177324
rect 184256 177284 184262 177296
rect 324406 177284 324412 177296
rect 324464 177284 324470 177336
rect 333238 177284 333244 177336
rect 333296 177324 333302 177336
rect 338114 177324 338120 177336
rect 333296 177296 338120 177324
rect 333296 177284 333302 177296
rect 338114 177284 338120 177296
rect 338172 177284 338178 177336
rect 134426 177012 134432 177064
rect 134484 177052 134490 177064
rect 165430 177052 165436 177064
rect 134484 177024 165436 177052
rect 134484 177012 134490 177024
rect 165430 177012 165436 177024
rect 165488 177012 165494 177064
rect 103330 176944 103336 176996
rect 103388 176984 103394 176996
rect 169202 176984 169208 176996
rect 103388 176956 169208 176984
rect 103388 176944 103394 176956
rect 169202 176944 169208 176956
rect 169260 176944 169266 176996
rect 108114 176876 108120 176928
rect 108172 176916 108178 176928
rect 184842 176916 184848 176928
rect 108172 176888 184848 176916
rect 108172 176876 108178 176888
rect 184842 176876 184848 176888
rect 184900 176876 184906 176928
rect 136082 176808 136088 176860
rect 136140 176848 136146 176860
rect 213914 176848 213920 176860
rect 136140 176820 213920 176848
rect 136140 176808 136146 176820
rect 213914 176808 213920 176820
rect 213972 176808 213978 176860
rect 125870 176740 125876 176792
rect 125928 176780 125934 176792
rect 214926 176780 214932 176792
rect 125928 176752 214932 176780
rect 125928 176740 125934 176752
rect 214926 176740 214932 176752
rect 214984 176740 214990 176792
rect 102042 176672 102048 176724
rect 102100 176712 102106 176724
rect 202230 176712 202236 176724
rect 102100 176684 202236 176712
rect 102100 176672 102106 176684
rect 202230 176672 202236 176684
rect 202288 176672 202294 176724
rect 132034 176264 132040 176316
rect 132092 176304 132098 176316
rect 165522 176304 165528 176316
rect 132092 176276 165528 176304
rect 132092 176264 132098 176276
rect 165522 176264 165528 176276
rect 165580 176264 165586 176316
rect 158898 176196 158904 176248
rect 158956 176236 158962 176248
rect 198090 176236 198096 176248
rect 158956 176208 198096 176236
rect 158956 176196 158962 176208
rect 198090 176196 198096 176208
rect 198148 176196 198154 176248
rect 238110 176196 238116 176248
rect 238168 176236 238174 176248
rect 249242 176236 249248 176248
rect 238168 176208 249248 176236
rect 238168 176196 238174 176208
rect 249242 176196 249248 176208
rect 249300 176196 249306 176248
rect 118418 176128 118424 176180
rect 118476 176168 118482 176180
rect 166258 176168 166264 176180
rect 118476 176140 166264 176168
rect 118476 176128 118482 176140
rect 166258 176128 166264 176140
rect 166316 176128 166322 176180
rect 239490 176128 239496 176180
rect 239548 176168 239554 176180
rect 249058 176168 249064 176180
rect 239548 176140 249064 176168
rect 239548 176128 239554 176140
rect 249058 176128 249064 176140
rect 249116 176128 249122 176180
rect 319438 176128 319444 176180
rect 319496 176168 319502 176180
rect 326154 176168 326160 176180
rect 319496 176140 326160 176168
rect 319496 176128 319502 176140
rect 326154 176128 326160 176140
rect 326212 176128 326218 176180
rect 121914 176060 121920 176112
rect 121972 176100 121978 176112
rect 170674 176100 170680 176112
rect 121972 176072 170680 176100
rect 121972 176060 121978 176072
rect 170674 176060 170680 176072
rect 170732 176060 170738 176112
rect 246390 176060 246396 176112
rect 246448 176100 246454 176112
rect 255590 176100 255596 176112
rect 246448 176072 255596 176100
rect 246448 176060 246454 176072
rect 255590 176060 255596 176072
rect 255648 176060 255654 176112
rect 312538 176060 312544 176112
rect 312596 176100 312602 176112
rect 321462 176100 321468 176112
rect 312596 176072 321468 176100
rect 312596 176060 312602 176072
rect 321462 176060 321468 176072
rect 321520 176060 321526 176112
rect 100754 175992 100760 176044
rect 100812 176032 100818 176044
rect 184198 176032 184204 176044
rect 100812 176004 184204 176032
rect 100812 175992 100818 176004
rect 184198 175992 184204 176004
rect 184256 175992 184262 176044
rect 184842 175992 184848 176044
rect 184900 176032 184906 176044
rect 214558 176032 214564 176044
rect 184900 176004 214564 176032
rect 184900 175992 184906 176004
rect 214558 175992 214564 176004
rect 214616 175992 214622 176044
rect 316678 175992 316684 176044
rect 316736 176032 316742 176044
rect 332870 176032 332876 176044
rect 316736 176004 332876 176032
rect 316736 175992 316742 176004
rect 332870 175992 332876 176004
rect 332928 175992 332934 176044
rect 11698 175924 11704 175976
rect 11756 175964 11762 175976
rect 111058 175964 111064 175976
rect 11756 175936 111064 175964
rect 11756 175924 11762 175936
rect 111058 175924 111064 175936
rect 111116 175924 111122 175976
rect 127066 175924 127072 175976
rect 127124 175964 127130 175976
rect 211890 175964 211896 175976
rect 127124 175936 211896 175964
rect 127124 175924 127130 175936
rect 211890 175924 211896 175936
rect 211948 175924 211954 175976
rect 236638 175924 236644 175976
rect 236696 175964 236702 175976
rect 256878 175964 256884 175976
rect 236696 175936 256884 175964
rect 236696 175924 236702 175936
rect 256878 175924 256884 175936
rect 256936 175924 256942 175976
rect 318058 175924 318064 175976
rect 318116 175964 318122 175976
rect 337010 175964 337016 175976
rect 318116 175936 337016 175964
rect 318116 175924 318122 175936
rect 337010 175924 337016 175936
rect 337068 175924 337074 175976
rect 165430 175176 165436 175228
rect 165488 175216 165494 175228
rect 213914 175216 213920 175228
rect 165488 175188 213920 175216
rect 165488 175176 165494 175188
rect 213914 175176 213920 175188
rect 213972 175176 213978 175228
rect 164878 175108 164884 175160
rect 164936 175148 164942 175160
rect 214006 175148 214012 175160
rect 164936 175120 214012 175148
rect 164936 175108 164942 175120
rect 214006 175108 214012 175120
rect 214064 175108 214070 175160
rect 291930 174020 291936 174072
rect 291988 174060 291994 174072
rect 307662 174060 307668 174072
rect 291988 174032 307668 174060
rect 291988 174020 291994 174032
rect 307662 174020 307668 174032
rect 307720 174020 307726 174072
rect 289170 173952 289176 174004
rect 289228 173992 289234 174004
rect 307478 173992 307484 174004
rect 289228 173964 307484 173992
rect 289228 173952 289234 173964
rect 307478 173952 307484 173964
rect 307536 173952 307542 174004
rect 269758 173884 269764 173936
rect 269816 173924 269822 173936
rect 307570 173924 307576 173936
rect 269816 173896 307576 173924
rect 269816 173884 269822 173896
rect 307570 173884 307576 173896
rect 307628 173884 307634 173936
rect 165522 173816 165528 173868
rect 165580 173856 165586 173868
rect 213914 173856 213920 173868
rect 165580 173828 213920 173856
rect 165580 173816 165586 173828
rect 213914 173816 213920 173828
rect 213972 173816 213978 173868
rect 252462 173816 252468 173868
rect 252520 173856 252526 173868
rect 263778 173856 263784 173868
rect 252520 173828 263784 173856
rect 252520 173816 252526 173828
rect 263778 173816 263784 173828
rect 263836 173816 263842 173868
rect 324314 173816 324320 173868
rect 324372 173856 324378 173868
rect 326154 173856 326160 173868
rect 324372 173828 326160 173856
rect 324372 173816 324378 173828
rect 326154 173816 326160 173828
rect 326212 173816 326218 173868
rect 295978 172660 295984 172712
rect 296036 172700 296042 172712
rect 307478 172700 307484 172712
rect 296036 172672 307484 172700
rect 296036 172660 296042 172672
rect 307478 172660 307484 172672
rect 307536 172660 307542 172712
rect 289078 172592 289084 172644
rect 289136 172632 289142 172644
rect 307570 172632 307576 172644
rect 289136 172604 307576 172632
rect 289136 172592 289142 172604
rect 307570 172592 307576 172604
rect 307628 172592 307634 172644
rect 266998 172524 267004 172576
rect 267056 172564 267062 172576
rect 307662 172564 307668 172576
rect 267056 172536 307668 172564
rect 267056 172524 267062 172536
rect 307662 172524 307668 172536
rect 307720 172524 307726 172576
rect 166534 172456 166540 172508
rect 166592 172496 166598 172508
rect 214006 172496 214012 172508
rect 166592 172468 214012 172496
rect 166592 172456 166598 172468
rect 214006 172456 214012 172468
rect 214064 172456 214070 172508
rect 177298 172388 177304 172440
rect 177356 172428 177362 172440
rect 213914 172428 213920 172440
rect 177356 172400 213920 172428
rect 177356 172388 177362 172400
rect 213914 172388 213920 172400
rect 213972 172388 213978 172440
rect 252462 172320 252468 172372
rect 252520 172360 252526 172372
rect 266354 172360 266360 172372
rect 252520 172332 266360 172360
rect 252520 172320 252526 172332
rect 266354 172320 266360 172332
rect 266412 172320 266418 172372
rect 296070 171232 296076 171284
rect 296128 171272 296134 171284
rect 306558 171272 306564 171284
rect 296128 171244 306564 171272
rect 296128 171232 296134 171244
rect 306558 171232 306564 171244
rect 306616 171232 306622 171284
rect 268378 171164 268384 171216
rect 268436 171204 268442 171216
rect 307570 171204 307576 171216
rect 268436 171176 307576 171204
rect 268436 171164 268442 171176
rect 307570 171164 307576 171176
rect 307628 171164 307634 171216
rect 264422 171096 264428 171148
rect 264480 171136 264486 171148
rect 307662 171136 307668 171148
rect 264480 171108 307668 171136
rect 264480 171096 264486 171108
rect 307662 171096 307668 171108
rect 307720 171096 307726 171148
rect 211890 171028 211896 171080
rect 211948 171068 211954 171080
rect 214466 171068 214472 171080
rect 211948 171040 214472 171068
rect 211948 171028 211954 171040
rect 214466 171028 214472 171040
rect 214524 171028 214530 171080
rect 252370 171028 252376 171080
rect 252428 171068 252434 171080
rect 265066 171068 265072 171080
rect 252428 171040 265072 171068
rect 252428 171028 252434 171040
rect 265066 171028 265072 171040
rect 265124 171028 265130 171080
rect 324314 171028 324320 171080
rect 324372 171068 324378 171080
rect 338114 171068 338120 171080
rect 324372 171040 338120 171068
rect 324372 171028 324378 171040
rect 338114 171028 338120 171040
rect 338172 171028 338178 171080
rect 252278 170824 252284 170876
rect 252336 170864 252342 170876
rect 256878 170864 256884 170876
rect 252336 170836 256884 170864
rect 252336 170824 252342 170836
rect 256878 170824 256884 170836
rect 256936 170824 256942 170876
rect 252462 170756 252468 170808
rect 252520 170796 252526 170808
rect 258258 170796 258264 170808
rect 252520 170768 258264 170796
rect 252520 170756 252526 170768
rect 258258 170756 258264 170768
rect 258316 170756 258322 170808
rect 300118 169872 300124 169924
rect 300176 169912 300182 169924
rect 307662 169912 307668 169924
rect 300176 169884 307668 169912
rect 300176 169872 300182 169884
rect 307662 169872 307668 169884
rect 307720 169872 307726 169924
rect 286410 169804 286416 169856
rect 286468 169844 286474 169856
rect 307294 169844 307300 169856
rect 286468 169816 307300 169844
rect 286468 169804 286474 169816
rect 307294 169804 307300 169816
rect 307352 169804 307358 169856
rect 259086 169736 259092 169788
rect 259144 169776 259150 169788
rect 262214 169776 262220 169788
rect 259144 169748 262220 169776
rect 259144 169736 259150 169748
rect 262214 169736 262220 169748
rect 262272 169736 262278 169788
rect 275370 169736 275376 169788
rect 275428 169776 275434 169788
rect 307478 169776 307484 169788
rect 275428 169748 307484 169776
rect 275428 169736 275434 169748
rect 307478 169736 307484 169748
rect 307536 169736 307542 169788
rect 166350 169668 166356 169720
rect 166408 169708 166414 169720
rect 214006 169708 214012 169720
rect 166408 169680 214012 169708
rect 166408 169668 166414 169680
rect 214006 169668 214012 169680
rect 214064 169668 214070 169720
rect 252370 169668 252376 169720
rect 252428 169708 252434 169720
rect 260834 169708 260840 169720
rect 252428 169680 260840 169708
rect 252428 169668 252434 169680
rect 260834 169668 260840 169680
rect 260892 169668 260898 169720
rect 324314 169668 324320 169720
rect 324372 169708 324378 169720
rect 345290 169708 345296 169720
rect 324372 169680 345296 169708
rect 324372 169668 324378 169680
rect 345290 169668 345296 169680
rect 345348 169668 345354 169720
rect 167914 169600 167920 169652
rect 167972 169640 167978 169652
rect 213914 169640 213920 169652
rect 167972 169612 213920 169640
rect 167972 169600 167978 169612
rect 213914 169600 213920 169612
rect 213972 169600 213978 169652
rect 252462 169056 252468 169108
rect 252520 169096 252526 169108
rect 258350 169096 258356 169108
rect 252520 169068 258356 169096
rect 252520 169056 252526 169068
rect 258350 169056 258356 169068
rect 258408 169056 258414 169108
rect 252462 168648 252468 168700
rect 252520 168688 252526 168700
rect 259730 168688 259736 168700
rect 252520 168660 259736 168688
rect 252520 168648 252526 168660
rect 259730 168648 259736 168660
rect 259788 168648 259794 168700
rect 290458 168512 290464 168564
rect 290516 168552 290522 168564
rect 307110 168552 307116 168564
rect 290516 168524 307116 168552
rect 290516 168512 290522 168524
rect 307110 168512 307116 168524
rect 307168 168512 307174 168564
rect 271322 168444 271328 168496
rect 271380 168484 271386 168496
rect 307662 168484 307668 168496
rect 271380 168456 307668 168484
rect 271380 168444 271386 168456
rect 307662 168444 307668 168456
rect 307720 168444 307726 168496
rect 262858 168376 262864 168428
rect 262916 168416 262922 168428
rect 307570 168416 307576 168428
rect 262916 168388 307576 168416
rect 262916 168376 262922 168388
rect 307570 168376 307576 168388
rect 307628 168376 307634 168428
rect 167730 168308 167736 168360
rect 167788 168348 167794 168360
rect 214006 168348 214012 168360
rect 167788 168320 214012 168348
rect 167788 168308 167794 168320
rect 214006 168308 214012 168320
rect 214064 168308 214070 168360
rect 252370 168308 252376 168360
rect 252428 168348 252434 168360
rect 263594 168348 263600 168360
rect 252428 168320 263600 168348
rect 252428 168308 252434 168320
rect 263594 168308 263600 168320
rect 263652 168308 263658 168360
rect 324314 168308 324320 168360
rect 324372 168348 324378 168360
rect 339586 168348 339592 168360
rect 324372 168320 339592 168348
rect 324372 168308 324378 168320
rect 339586 168308 339592 168320
rect 339644 168308 339650 168360
rect 170674 168240 170680 168292
rect 170732 168280 170738 168292
rect 213914 168280 213920 168292
rect 170732 168252 213920 168280
rect 170732 168240 170738 168252
rect 213914 168240 213920 168252
rect 213972 168240 213978 168292
rect 252462 168240 252468 168292
rect 252520 168280 252526 168292
rect 262398 168280 262404 168292
rect 252520 168252 262404 168280
rect 252520 168240 252526 168252
rect 262398 168240 262404 168252
rect 262456 168240 262462 168292
rect 324406 168240 324412 168292
rect 324464 168280 324470 168292
rect 331214 168280 331220 168292
rect 324464 168252 331220 168280
rect 324464 168240 324470 168252
rect 331214 168240 331220 168252
rect 331272 168240 331278 168292
rect 252462 167220 252468 167272
rect 252520 167260 252526 167272
rect 259086 167260 259092 167272
rect 252520 167232 259092 167260
rect 252520 167220 252526 167232
rect 259086 167220 259092 167232
rect 259144 167220 259150 167272
rect 283742 167152 283748 167204
rect 283800 167192 283806 167204
rect 307478 167192 307484 167204
rect 283800 167164 307484 167192
rect 283800 167152 283806 167164
rect 307478 167152 307484 167164
rect 307536 167152 307542 167204
rect 281074 167084 281080 167136
rect 281132 167124 281138 167136
rect 307662 167124 307668 167136
rect 281132 167096 307668 167124
rect 281132 167084 281138 167096
rect 307662 167084 307668 167096
rect 307720 167084 307726 167136
rect 276658 167016 276664 167068
rect 276716 167056 276722 167068
rect 307294 167056 307300 167068
rect 276716 167028 307300 167056
rect 276716 167016 276722 167028
rect 307294 167016 307300 167028
rect 307352 167016 307358 167068
rect 166258 166948 166264 167000
rect 166316 166988 166322 167000
rect 214006 166988 214012 167000
rect 166316 166960 214012 166988
rect 166316 166948 166322 166960
rect 214006 166948 214012 166960
rect 214064 166948 214070 167000
rect 252370 166948 252376 167000
rect 252428 166988 252434 167000
rect 261018 166988 261024 167000
rect 252428 166960 261024 166988
rect 252428 166948 252434 166960
rect 261018 166948 261024 166960
rect 261076 166948 261082 167000
rect 324314 166948 324320 167000
rect 324372 166988 324378 167000
rect 346670 166988 346676 167000
rect 324372 166960 346676 166988
rect 324372 166948 324378 166960
rect 346670 166948 346676 166960
rect 346728 166948 346734 167000
rect 464338 166948 464344 167000
rect 464396 166988 464402 167000
rect 580166 166988 580172 167000
rect 464396 166960 580172 166988
rect 464396 166948 464402 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 170582 166880 170588 166932
rect 170640 166920 170646 166932
rect 213914 166920 213920 166932
rect 170640 166892 213920 166920
rect 170640 166880 170646 166892
rect 213914 166880 213920 166892
rect 213972 166880 213978 166932
rect 252462 166812 252468 166864
rect 252520 166852 252526 166864
rect 259454 166852 259460 166864
rect 252520 166824 259460 166852
rect 252520 166812 252526 166824
rect 259454 166812 259460 166824
rect 259512 166812 259518 166864
rect 302878 165724 302884 165776
rect 302936 165764 302942 165776
rect 307110 165764 307116 165776
rect 302936 165736 307116 165764
rect 302936 165724 302942 165736
rect 307110 165724 307116 165736
rect 307168 165724 307174 165776
rect 278222 165656 278228 165708
rect 278280 165696 278286 165708
rect 307570 165696 307576 165708
rect 278280 165668 307576 165696
rect 278280 165656 278286 165668
rect 307570 165656 307576 165668
rect 307628 165656 307634 165708
rect 260190 165588 260196 165640
rect 260248 165628 260254 165640
rect 307662 165628 307668 165640
rect 260248 165600 307668 165628
rect 260248 165588 260254 165600
rect 307662 165588 307668 165600
rect 307720 165588 307726 165640
rect 166442 165520 166448 165572
rect 166500 165560 166506 165572
rect 213914 165560 213920 165572
rect 166500 165532 213920 165560
rect 166500 165520 166506 165532
rect 213914 165520 213920 165532
rect 213972 165520 213978 165572
rect 252370 165520 252376 165572
rect 252428 165560 252434 165572
rect 270494 165560 270500 165572
rect 252428 165532 270500 165560
rect 252428 165520 252434 165532
rect 270494 165520 270500 165532
rect 270552 165520 270558 165572
rect 324406 165520 324412 165572
rect 324464 165560 324470 165572
rect 346578 165560 346584 165572
rect 324464 165532 346584 165560
rect 324464 165520 324470 165532
rect 346578 165520 346584 165532
rect 346636 165520 346642 165572
rect 169294 165452 169300 165504
rect 169352 165492 169358 165504
rect 214006 165492 214012 165504
rect 169352 165464 214012 165492
rect 169352 165452 169358 165464
rect 214006 165452 214012 165464
rect 214064 165452 214070 165504
rect 252462 165452 252468 165504
rect 252520 165492 252526 165504
rect 261110 165492 261116 165504
rect 252520 165464 261116 165492
rect 252520 165452 252526 165464
rect 261110 165452 261116 165464
rect 261168 165452 261174 165504
rect 324314 165452 324320 165504
rect 324372 165492 324378 165504
rect 343910 165492 343916 165504
rect 324372 165464 343916 165492
rect 324372 165452 324378 165464
rect 343910 165452 343916 165464
rect 343968 165452 343974 165504
rect 251358 165384 251364 165436
rect 251416 165424 251422 165436
rect 254118 165424 254124 165436
rect 251416 165396 254124 165424
rect 251416 165384 251422 165396
rect 254118 165384 254124 165396
rect 254176 165384 254182 165436
rect 269850 164840 269856 164892
rect 269908 164880 269914 164892
rect 307386 164880 307392 164892
rect 269908 164852 307392 164880
rect 269908 164840 269914 164852
rect 307386 164840 307392 164852
rect 307444 164840 307450 164892
rect 305730 164296 305736 164348
rect 305788 164336 305794 164348
rect 307110 164336 307116 164348
rect 305788 164308 307116 164336
rect 305788 164296 305794 164308
rect 307110 164296 307116 164308
rect 307168 164296 307174 164348
rect 287974 164228 287980 164280
rect 288032 164268 288038 164280
rect 307662 164268 307668 164280
rect 288032 164240 307668 164268
rect 288032 164228 288038 164240
rect 307662 164228 307668 164240
rect 307720 164228 307726 164280
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 14458 164200 14464 164212
rect 3292 164172 14464 164200
rect 3292 164160 3298 164172
rect 14458 164160 14464 164172
rect 14516 164160 14522 164212
rect 170490 164160 170496 164212
rect 170548 164200 170554 164212
rect 213914 164200 213920 164212
rect 170548 164172 213920 164200
rect 170548 164160 170554 164172
rect 213914 164160 213920 164172
rect 213972 164160 213978 164212
rect 252370 164160 252376 164212
rect 252428 164200 252434 164212
rect 266538 164200 266544 164212
rect 252428 164172 266544 164200
rect 252428 164160 252434 164172
rect 266538 164160 266544 164172
rect 266596 164160 266602 164212
rect 324406 164160 324412 164212
rect 324464 164200 324470 164212
rect 336918 164200 336924 164212
rect 324464 164172 336924 164200
rect 324464 164160 324470 164172
rect 336918 164160 336924 164172
rect 336976 164160 336982 164212
rect 252278 164092 252284 164144
rect 252336 164132 252342 164144
rect 265250 164132 265256 164144
rect 252336 164104 265256 164132
rect 252336 164092 252342 164104
rect 265250 164092 265256 164104
rect 265308 164092 265314 164144
rect 324314 164092 324320 164144
rect 324372 164132 324378 164144
rect 332870 164132 332876 164144
rect 324372 164104 332876 164132
rect 324372 164092 324378 164104
rect 332870 164092 332876 164104
rect 332928 164092 332934 164144
rect 252462 164024 252468 164076
rect 252520 164064 252526 164076
rect 263870 164064 263876 164076
rect 252520 164036 263876 164064
rect 252520 164024 252526 164036
rect 263870 164024 263876 164036
rect 263928 164024 263934 164076
rect 301498 163004 301504 163056
rect 301556 163044 301562 163056
rect 307570 163044 307576 163056
rect 301556 163016 307576 163044
rect 301556 163004 301562 163016
rect 307570 163004 307576 163016
rect 307628 163004 307634 163056
rect 271230 162936 271236 162988
rect 271288 162976 271294 162988
rect 306742 162976 306748 162988
rect 271288 162948 306748 162976
rect 271288 162936 271294 162948
rect 306742 162936 306748 162948
rect 306800 162936 306806 162988
rect 257522 162868 257528 162920
rect 257580 162908 257586 162920
rect 307662 162908 307668 162920
rect 257580 162880 307668 162908
rect 257580 162868 257586 162880
rect 307662 162868 307668 162880
rect 307720 162868 307726 162920
rect 167638 162800 167644 162852
rect 167696 162840 167702 162852
rect 213914 162840 213920 162852
rect 167696 162812 213920 162840
rect 167696 162800 167702 162812
rect 213914 162800 213920 162812
rect 213972 162800 213978 162852
rect 324406 162800 324412 162852
rect 324464 162840 324470 162852
rect 335538 162840 335544 162852
rect 324464 162812 335544 162840
rect 324464 162800 324470 162812
rect 335538 162800 335544 162812
rect 335596 162800 335602 162852
rect 170398 162732 170404 162784
rect 170456 162772 170462 162784
rect 214006 162772 214012 162784
rect 170456 162744 214012 162772
rect 170456 162732 170462 162744
rect 214006 162732 214012 162744
rect 214064 162732 214070 162784
rect 252462 162732 252468 162784
rect 252520 162772 252526 162784
rect 267734 162772 267740 162784
rect 252520 162744 267740 162772
rect 252520 162732 252526 162744
rect 267734 162732 267740 162744
rect 267792 162732 267798 162784
rect 324314 162732 324320 162784
rect 324372 162772 324378 162784
rect 330110 162772 330116 162784
rect 324372 162744 330116 162772
rect 324372 162732 324378 162744
rect 330110 162732 330116 162744
rect 330168 162732 330174 162784
rect 297450 161576 297456 161628
rect 297508 161616 297514 161628
rect 307478 161616 307484 161628
rect 297508 161588 307484 161616
rect 297508 161576 297514 161588
rect 307478 161576 307484 161588
rect 307536 161576 307542 161628
rect 264238 161508 264244 161560
rect 264296 161548 264302 161560
rect 307570 161548 307576 161560
rect 264296 161520 307576 161548
rect 264296 161508 264302 161520
rect 307570 161508 307576 161520
rect 307628 161508 307634 161560
rect 258902 161440 258908 161492
rect 258960 161480 258966 161492
rect 307662 161480 307668 161492
rect 258960 161452 307668 161480
rect 258960 161440 258966 161452
rect 307662 161440 307668 161452
rect 307720 161440 307726 161492
rect 188430 161372 188436 161424
rect 188488 161412 188494 161424
rect 213914 161412 213920 161424
rect 188488 161384 213920 161412
rect 188488 161372 188494 161384
rect 213914 161372 213920 161384
rect 213972 161372 213978 161424
rect 252370 161372 252376 161424
rect 252428 161412 252434 161424
rect 270678 161412 270684 161424
rect 252428 161384 270684 161412
rect 252428 161372 252434 161384
rect 270678 161372 270684 161384
rect 270736 161372 270742 161424
rect 324314 161372 324320 161424
rect 324372 161412 324378 161424
rect 337010 161412 337016 161424
rect 324372 161384 337016 161412
rect 324372 161372 324378 161384
rect 337010 161372 337016 161384
rect 337068 161372 337074 161424
rect 324406 161304 324412 161356
rect 324464 161344 324470 161356
rect 332778 161344 332784 161356
rect 324464 161316 332784 161344
rect 324464 161304 324470 161316
rect 332778 161304 332784 161316
rect 332836 161304 332842 161356
rect 252002 160964 252008 161016
rect 252060 161004 252066 161016
rect 255314 161004 255320 161016
rect 252060 160976 255320 161004
rect 252060 160964 252066 160976
rect 255314 160964 255320 160976
rect 255372 160964 255378 161016
rect 252462 160760 252468 160812
rect 252520 160800 252526 160812
rect 258166 160800 258172 160812
rect 252520 160772 258172 160800
rect 252520 160760 252526 160772
rect 258166 160760 258172 160772
rect 258224 160760 258230 160812
rect 167822 160692 167828 160744
rect 167880 160732 167886 160744
rect 214650 160732 214656 160744
rect 167880 160704 214656 160732
rect 167880 160692 167886 160704
rect 214650 160692 214656 160704
rect 214708 160692 214714 160744
rect 291838 160216 291844 160268
rect 291896 160256 291902 160268
rect 307662 160256 307668 160268
rect 291896 160228 307668 160256
rect 291896 160216 291902 160228
rect 307662 160216 307668 160228
rect 307720 160216 307726 160268
rect 265618 160148 265624 160200
rect 265676 160188 265682 160200
rect 306558 160188 306564 160200
rect 265676 160160 306564 160188
rect 265676 160148 265682 160160
rect 306558 160148 306564 160160
rect 306616 160148 306622 160200
rect 258718 160080 258724 160132
rect 258776 160120 258782 160132
rect 307570 160120 307576 160132
rect 258776 160092 307576 160120
rect 258776 160080 258782 160092
rect 307570 160080 307576 160092
rect 307628 160080 307634 160132
rect 173250 160012 173256 160064
rect 173308 160052 173314 160064
rect 213914 160052 213920 160064
rect 173308 160024 213920 160052
rect 173308 160012 173314 160024
rect 213914 160012 213920 160024
rect 213972 160012 213978 160064
rect 252462 160012 252468 160064
rect 252520 160052 252526 160064
rect 274818 160052 274824 160064
rect 252520 160024 274824 160052
rect 252520 160012 252526 160024
rect 274818 160012 274824 160024
rect 274876 160012 274882 160064
rect 298830 159332 298836 159384
rect 298888 159372 298894 159384
rect 307202 159372 307208 159384
rect 298888 159344 307208 159372
rect 298888 159332 298894 159344
rect 307202 159332 307208 159344
rect 307260 159332 307266 159384
rect 262950 158788 262956 158840
rect 263008 158828 263014 158840
rect 307570 158828 307576 158840
rect 263008 158800 307576 158828
rect 263008 158788 263014 158800
rect 307570 158788 307576 158800
rect 307628 158788 307634 158840
rect 254578 158720 254584 158772
rect 254636 158760 254642 158772
rect 307662 158760 307668 158772
rect 254636 158732 307668 158760
rect 254636 158720 254642 158732
rect 307662 158720 307668 158732
rect 307720 158720 307726 158772
rect 169202 158652 169208 158704
rect 169260 158692 169266 158704
rect 213914 158692 213920 158704
rect 169260 158664 213920 158692
rect 169260 158652 169266 158664
rect 213914 158652 213920 158664
rect 213972 158652 213978 158704
rect 252462 158652 252468 158704
rect 252520 158692 252526 158704
rect 276198 158692 276204 158704
rect 252520 158664 276204 158692
rect 252520 158652 252526 158664
rect 276198 158652 276204 158664
rect 276256 158652 276262 158704
rect 324406 158652 324412 158704
rect 324464 158692 324470 158704
rect 350626 158692 350632 158704
rect 324464 158664 350632 158692
rect 324464 158652 324470 158664
rect 350626 158652 350632 158664
rect 350684 158652 350690 158704
rect 202230 158584 202236 158636
rect 202288 158624 202294 158636
rect 214006 158624 214012 158636
rect 202288 158596 214012 158624
rect 202288 158584 202294 158596
rect 214006 158584 214012 158596
rect 214064 158584 214070 158636
rect 324314 158584 324320 158636
rect 324372 158624 324378 158636
rect 334066 158624 334072 158636
rect 324372 158596 334072 158624
rect 324372 158584 324378 158596
rect 334066 158584 334072 158596
rect 334124 158584 334130 158636
rect 293402 157496 293408 157548
rect 293460 157536 293466 157548
rect 307662 157536 307668 157548
rect 293460 157508 307668 157536
rect 293460 157496 293466 157508
rect 307662 157496 307668 157508
rect 307720 157496 307726 157548
rect 264330 157428 264336 157480
rect 264388 157468 264394 157480
rect 306926 157468 306932 157480
rect 264388 157440 306932 157468
rect 264388 157428 264394 157440
rect 306926 157428 306932 157440
rect 306984 157428 306990 157480
rect 258810 157360 258816 157412
rect 258868 157400 258874 157412
rect 307570 157400 307576 157412
rect 258868 157372 307576 157400
rect 258868 157360 258874 157372
rect 307570 157360 307576 157372
rect 307628 157360 307634 157412
rect 169110 157292 169116 157344
rect 169168 157332 169174 157344
rect 214006 157332 214012 157344
rect 169168 157304 214012 157332
rect 169168 157292 169174 157304
rect 214006 157292 214012 157304
rect 214064 157292 214070 157344
rect 252370 157292 252376 157344
rect 252428 157332 252434 157344
rect 272058 157332 272064 157344
rect 252428 157304 272064 157332
rect 252428 157292 252434 157304
rect 272058 157292 272064 157304
rect 272116 157292 272122 157344
rect 184198 157224 184204 157276
rect 184256 157264 184262 157276
rect 213914 157264 213920 157276
rect 184256 157236 213920 157264
rect 184256 157224 184262 157236
rect 213914 157224 213920 157236
rect 213972 157224 213978 157276
rect 252462 157224 252468 157276
rect 252520 157264 252526 157276
rect 265158 157264 265164 157276
rect 252520 157236 265164 157264
rect 252520 157224 252526 157236
rect 265158 157224 265164 157236
rect 265216 157224 265222 157276
rect 324314 157224 324320 157276
rect 324372 157264 324378 157276
rect 349338 157264 349344 157276
rect 324372 157236 349344 157264
rect 324372 157224 324378 157236
rect 349338 157224 349344 157236
rect 349396 157224 349402 157276
rect 324314 156816 324320 156868
rect 324372 156856 324378 156868
rect 325970 156856 325976 156868
rect 324372 156828 325976 156856
rect 324372 156816 324378 156828
rect 325970 156816 325976 156828
rect 326028 156816 326034 156868
rect 300762 156068 300768 156120
rect 300820 156108 300826 156120
rect 307662 156108 307668 156120
rect 300820 156080 307668 156108
rect 300820 156068 300826 156080
rect 307662 156068 307668 156080
rect 307720 156068 307726 156120
rect 268470 156000 268476 156052
rect 268528 156040 268534 156052
rect 307478 156040 307484 156052
rect 268528 156012 307484 156040
rect 268528 156000 268534 156012
rect 307478 156000 307484 156012
rect 307536 156000 307542 156052
rect 260098 155932 260104 155984
rect 260156 155972 260162 155984
rect 307570 155972 307576 155984
rect 260156 155944 307576 155972
rect 260156 155932 260162 155944
rect 307570 155932 307576 155944
rect 307628 155932 307634 155984
rect 171778 155864 171784 155916
rect 171836 155904 171842 155916
rect 213914 155904 213920 155916
rect 171836 155876 213920 155904
rect 171836 155864 171842 155876
rect 213914 155864 213920 155876
rect 213972 155864 213978 155916
rect 252462 155864 252468 155916
rect 252520 155904 252526 155916
rect 254026 155904 254032 155916
rect 252520 155876 254032 155904
rect 252520 155864 252526 155876
rect 254026 155864 254032 155876
rect 254084 155864 254090 155916
rect 324406 155864 324412 155916
rect 324464 155904 324470 155916
rect 341150 155904 341156 155916
rect 324464 155876 341156 155904
rect 324464 155864 324470 155876
rect 341150 155864 341156 155876
rect 341208 155864 341214 155916
rect 251542 155796 251548 155848
rect 251600 155836 251606 155848
rect 254210 155836 254216 155848
rect 251600 155808 254216 155836
rect 251600 155796 251606 155808
rect 254210 155796 254216 155808
rect 254268 155796 254274 155848
rect 324314 155796 324320 155848
rect 324372 155836 324378 155848
rect 339770 155836 339776 155848
rect 324372 155808 339776 155836
rect 324372 155796 324378 155808
rect 339770 155796 339776 155808
rect 339828 155796 339834 155848
rect 252462 155728 252468 155780
rect 252520 155768 252526 155780
rect 266446 155768 266452 155780
rect 252520 155740 266452 155768
rect 252520 155728 252526 155740
rect 266446 155728 266452 155740
rect 266504 155728 266510 155780
rect 282454 155184 282460 155236
rect 282512 155224 282518 155236
rect 307386 155224 307392 155236
rect 282512 155196 307392 155224
rect 282512 155184 282518 155196
rect 307386 155184 307392 155196
rect 307444 155184 307450 155236
rect 267090 154640 267096 154692
rect 267148 154680 267154 154692
rect 306558 154680 306564 154692
rect 267148 154652 306564 154680
rect 267148 154640 267154 154652
rect 306558 154640 306564 154652
rect 306616 154640 306622 154692
rect 254854 154572 254860 154624
rect 254912 154612 254918 154624
rect 307662 154612 307668 154624
rect 254912 154584 307668 154612
rect 254912 154572 254918 154584
rect 307662 154572 307668 154584
rect 307720 154572 307726 154624
rect 324314 154504 324320 154556
rect 324372 154544 324378 154556
rect 353386 154544 353392 154556
rect 324372 154516 353392 154544
rect 324372 154504 324378 154516
rect 353386 154504 353392 154516
rect 353444 154504 353450 154556
rect 252462 154436 252468 154488
rect 252520 154476 252526 154488
rect 269206 154476 269212 154488
rect 252520 154448 269212 154476
rect 252520 154436 252526 154448
rect 269206 154436 269212 154448
rect 269264 154436 269270 154488
rect 251818 153824 251824 153876
rect 251876 153864 251882 153876
rect 300762 153864 300768 153876
rect 251876 153836 300768 153864
rect 251876 153824 251882 153836
rect 300762 153824 300768 153836
rect 300820 153824 300826 153876
rect 324314 153416 324320 153468
rect 324372 153456 324378 153468
rect 327350 153456 327356 153468
rect 324372 153428 327356 153456
rect 324372 153416 324378 153428
rect 327350 153416 327356 153428
rect 327408 153416 327414 153468
rect 300394 153348 300400 153400
rect 300452 153388 300458 153400
rect 307570 153388 307576 153400
rect 300452 153360 307576 153388
rect 300452 153348 300458 153360
rect 307570 153348 307576 153360
rect 307628 153348 307634 153400
rect 178862 153280 178868 153332
rect 178920 153320 178926 153332
rect 214006 153320 214012 153332
rect 178920 153292 214012 153320
rect 178920 153280 178926 153292
rect 214006 153280 214012 153292
rect 214064 153280 214070 153332
rect 297634 153280 297640 153332
rect 297692 153320 297698 153332
rect 307662 153320 307668 153332
rect 297692 153292 307668 153320
rect 297692 153280 297698 153292
rect 307662 153280 307668 153292
rect 307720 153280 307726 153332
rect 175918 153212 175924 153264
rect 175976 153252 175982 153264
rect 213914 153252 213920 153264
rect 175976 153224 213920 153252
rect 175976 153212 175982 153224
rect 213914 153212 213920 153224
rect 213972 153212 213978 153264
rect 254762 153212 254768 153264
rect 254820 153252 254826 153264
rect 306558 153252 306564 153264
rect 254820 153224 306564 153252
rect 254820 153212 254826 153224
rect 306558 153212 306564 153224
rect 306616 153212 306622 153264
rect 252370 153144 252376 153196
rect 252428 153184 252434 153196
rect 273530 153184 273536 153196
rect 252428 153156 273536 153184
rect 252428 153144 252434 153156
rect 273530 153144 273536 153156
rect 273588 153144 273594 153196
rect 324406 153144 324412 153196
rect 324464 153184 324470 153196
rect 350718 153184 350724 153196
rect 324464 153156 350724 153184
rect 324464 153144 324470 153156
rect 350718 153144 350724 153156
rect 350776 153144 350782 153196
rect 252462 153076 252468 153128
rect 252520 153116 252526 153128
rect 267918 153116 267924 153128
rect 252520 153088 267924 153116
rect 252520 153076 252526 153088
rect 267918 153076 267924 153088
rect 267976 153076 267982 153128
rect 296162 151920 296168 151972
rect 296220 151960 296226 151972
rect 306558 151960 306564 151972
rect 296220 151932 306564 151960
rect 296220 151920 296226 151932
rect 306558 151920 306564 151932
rect 306616 151920 306622 151972
rect 184290 151852 184296 151904
rect 184348 151892 184354 151904
rect 213914 151892 213920 151904
rect 184348 151864 213920 151892
rect 184348 151852 184354 151864
rect 213914 151852 213920 151864
rect 213972 151852 213978 151904
rect 272794 151852 272800 151904
rect 272852 151892 272858 151904
rect 307662 151892 307668 151904
rect 272852 151864 307668 151892
rect 272852 151852 272858 151864
rect 307662 151852 307668 151864
rect 307720 151852 307726 151904
rect 177298 151784 177304 151836
rect 177356 151824 177362 151836
rect 214006 151824 214012 151836
rect 177356 151796 214012 151824
rect 177356 151784 177362 151796
rect 214006 151784 214012 151796
rect 214064 151784 214070 151836
rect 256142 151784 256148 151836
rect 256200 151824 256206 151836
rect 307478 151824 307484 151836
rect 256200 151796 307484 151824
rect 256200 151784 256206 151796
rect 307478 151784 307484 151796
rect 307536 151784 307542 151836
rect 252462 151716 252468 151768
rect 252520 151756 252526 151768
rect 281626 151756 281632 151768
rect 252520 151728 281632 151756
rect 252520 151716 252526 151728
rect 281626 151716 281632 151728
rect 281684 151716 281690 151768
rect 324314 151716 324320 151768
rect 324372 151756 324378 151768
rect 328638 151756 328644 151768
rect 324372 151728 328644 151756
rect 324372 151716 324378 151728
rect 328638 151716 328644 151728
rect 328696 151716 328702 151768
rect 252370 151648 252376 151700
rect 252428 151688 252434 151700
rect 255406 151688 255412 151700
rect 252428 151660 255412 151688
rect 252428 151648 252434 151660
rect 255406 151648 255412 151660
rect 255464 151648 255470 151700
rect 251358 151444 251364 151496
rect 251416 151484 251422 151496
rect 253934 151484 253940 151496
rect 251416 151456 253940 151484
rect 251416 151444 251422 151456
rect 253934 151444 253940 151456
rect 253992 151444 253998 151496
rect 300302 150560 300308 150612
rect 300360 150600 300366 150612
rect 307662 150600 307668 150612
rect 300360 150572 307668 150600
rect 300360 150560 300366 150572
rect 307662 150560 307668 150572
rect 307720 150560 307726 150612
rect 273990 150492 273996 150544
rect 274048 150532 274054 150544
rect 307478 150532 307484 150544
rect 274048 150504 307484 150532
rect 274048 150492 274054 150504
rect 307478 150492 307484 150504
rect 307536 150492 307542 150544
rect 199562 150424 199568 150476
rect 199620 150464 199626 150476
rect 213914 150464 213920 150476
rect 199620 150436 213920 150464
rect 199620 150424 199626 150436
rect 213914 150424 213920 150436
rect 213972 150424 213978 150476
rect 256050 150424 256056 150476
rect 256108 150464 256114 150476
rect 307570 150464 307576 150476
rect 256108 150436 307576 150464
rect 256108 150424 256114 150436
rect 307570 150424 307576 150436
rect 307628 150424 307634 150476
rect 3510 150356 3516 150408
rect 3568 150396 3574 150408
rect 21358 150396 21364 150408
rect 3568 150368 21364 150396
rect 3568 150356 3574 150368
rect 21358 150356 21364 150368
rect 21416 150356 21422 150408
rect 181438 150356 181444 150408
rect 181496 150396 181502 150408
rect 214006 150396 214012 150408
rect 181496 150368 214012 150396
rect 181496 150356 181502 150368
rect 214006 150356 214012 150368
rect 214064 150356 214070 150408
rect 252462 150356 252468 150408
rect 252520 150396 252526 150408
rect 277486 150396 277492 150408
rect 252520 150368 277492 150396
rect 252520 150356 252526 150368
rect 277486 150356 277492 150368
rect 277544 150356 277550 150408
rect 324314 150356 324320 150408
rect 324372 150396 324378 150408
rect 334250 150396 334256 150408
rect 324372 150368 334256 150396
rect 324372 150356 324378 150368
rect 334250 150356 334256 150368
rect 334308 150356 334314 150408
rect 252094 150288 252100 150340
rect 252152 150328 252158 150340
rect 255498 150328 255504 150340
rect 252152 150300 255504 150328
rect 252152 150288 252158 150300
rect 255498 150288 255504 150300
rect 255556 150288 255562 150340
rect 324406 150288 324412 150340
rect 324464 150328 324470 150340
rect 331306 150328 331312 150340
rect 324464 150300 331312 150328
rect 324464 150288 324470 150300
rect 331306 150288 331312 150300
rect 331364 150288 331370 150340
rect 252278 150220 252284 150272
rect 252336 150260 252342 150272
rect 255590 150260 255596 150272
rect 252336 150232 255596 150260
rect 252336 150220 252342 150232
rect 255590 150220 255596 150232
rect 255648 150220 255654 150272
rect 275462 149676 275468 149728
rect 275520 149716 275526 149728
rect 307202 149716 307208 149728
rect 275520 149688 307208 149716
rect 275520 149676 275526 149688
rect 307202 149676 307208 149688
rect 307260 149676 307266 149728
rect 255314 149336 255320 149388
rect 255372 149376 255378 149388
rect 258074 149376 258080 149388
rect 255372 149348 258080 149376
rect 255372 149336 255378 149348
rect 258074 149336 258080 149348
rect 258132 149336 258138 149388
rect 297726 149132 297732 149184
rect 297784 149172 297790 149184
rect 307478 149172 307484 149184
rect 297784 149144 307484 149172
rect 297784 149132 297790 149144
rect 307478 149132 307484 149144
rect 307536 149132 307542 149184
rect 254670 149064 254676 149116
rect 254728 149104 254734 149116
rect 306558 149104 306564 149116
rect 254728 149076 306564 149104
rect 254728 149064 254734 149076
rect 306558 149064 306564 149076
rect 306616 149064 306622 149116
rect 198090 148996 198096 149048
rect 198148 149036 198154 149048
rect 213914 149036 213920 149048
rect 198148 149008 213920 149036
rect 198148 148996 198154 149008
rect 213914 148996 213920 149008
rect 213972 148996 213978 149048
rect 252370 148996 252376 149048
rect 252428 149036 252434 149048
rect 280246 149036 280252 149048
rect 252428 149008 280252 149036
rect 252428 148996 252434 149008
rect 280246 148996 280252 149008
rect 280304 148996 280310 149048
rect 252462 148928 252468 148980
rect 252520 148968 252526 148980
rect 278866 148968 278872 148980
rect 252520 148940 278872 148968
rect 252520 148928 252526 148940
rect 278866 148928 278872 148940
rect 278924 148928 278930 148980
rect 324314 148928 324320 148980
rect 324372 148968 324378 148980
rect 347958 148968 347964 148980
rect 324372 148940 347964 148968
rect 324372 148928 324378 148940
rect 347958 148928 347964 148940
rect 348016 148928 348022 148980
rect 252278 148860 252284 148912
rect 252336 148900 252342 148912
rect 256786 148900 256792 148912
rect 252336 148872 256792 148900
rect 252336 148860 252342 148872
rect 256786 148860 256792 148872
rect 256844 148860 256850 148912
rect 258994 148316 259000 148368
rect 259052 148356 259058 148368
rect 306650 148356 306656 148368
rect 259052 148328 306656 148356
rect 259052 148316 259058 148328
rect 306650 148316 306656 148328
rect 306708 148316 306714 148368
rect 257338 147772 257344 147824
rect 257396 147812 257402 147824
rect 307662 147812 307668 147824
rect 257396 147784 307668 147812
rect 257396 147772 257402 147784
rect 307662 147772 307668 147784
rect 307720 147772 307726 147824
rect 167638 147636 167644 147688
rect 167696 147676 167702 147688
rect 213914 147676 213920 147688
rect 167696 147648 213920 147676
rect 167696 147636 167702 147648
rect 213914 147636 213920 147648
rect 213972 147636 213978 147688
rect 304350 147636 304356 147688
rect 304408 147676 304414 147688
rect 307294 147676 307300 147688
rect 304408 147648 307300 147676
rect 304408 147636 304414 147648
rect 307294 147636 307300 147648
rect 307352 147636 307358 147688
rect 324314 147568 324320 147620
rect 324372 147608 324378 147620
rect 335354 147608 335360 147620
rect 324372 147580 335360 147608
rect 324372 147568 324378 147580
rect 335354 147568 335360 147580
rect 335412 147568 335418 147620
rect 252462 147500 252468 147552
rect 252520 147540 252526 147552
rect 273346 147540 273352 147552
rect 252520 147512 273352 147540
rect 252520 147500 252526 147512
rect 273346 147500 273352 147512
rect 273404 147500 273410 147552
rect 252186 146888 252192 146940
rect 252244 146928 252250 146940
rect 260926 146928 260932 146940
rect 252244 146900 260932 146928
rect 252244 146888 252250 146900
rect 260926 146888 260932 146900
rect 260984 146888 260990 146940
rect 301774 146616 301780 146668
rect 301832 146656 301838 146668
rect 307570 146656 307576 146668
rect 301832 146628 307576 146656
rect 301832 146616 301838 146628
rect 307570 146616 307576 146628
rect 307628 146616 307634 146668
rect 210602 146344 210608 146396
rect 210660 146384 210666 146396
rect 214006 146384 214012 146396
rect 210660 146356 214012 146384
rect 210660 146344 210666 146356
rect 214006 146344 214012 146356
rect 214064 146344 214070 146396
rect 261478 146344 261484 146396
rect 261536 146384 261542 146396
rect 307294 146384 307300 146396
rect 261536 146356 307300 146384
rect 261536 146344 261542 146356
rect 307294 146344 307300 146356
rect 307352 146344 307358 146396
rect 174538 146276 174544 146328
rect 174596 146316 174602 146328
rect 213914 146316 213920 146328
rect 174596 146288 213920 146316
rect 174596 146276 174602 146288
rect 213914 146276 213920 146288
rect 213972 146276 213978 146328
rect 256234 146276 256240 146328
rect 256292 146316 256298 146328
rect 306926 146316 306932 146328
rect 256292 146288 306932 146316
rect 256292 146276 256298 146288
rect 306926 146276 306932 146288
rect 306984 146276 306990 146328
rect 252462 146208 252468 146260
rect 252520 146248 252526 146260
rect 280154 146248 280160 146260
rect 252520 146220 280160 146248
rect 252520 146208 252526 146220
rect 280154 146208 280160 146220
rect 280212 146208 280218 146260
rect 324314 146208 324320 146260
rect 324372 146248 324378 146260
rect 342346 146248 342352 146260
rect 324372 146220 342352 146248
rect 324372 146208 324378 146220
rect 342346 146208 342352 146220
rect 342404 146208 342410 146260
rect 252370 146140 252376 146192
rect 252428 146180 252434 146192
rect 270586 146180 270592 146192
rect 252428 146152 270592 146180
rect 252428 146140 252434 146152
rect 270586 146140 270592 146152
rect 270644 146140 270650 146192
rect 252278 146072 252284 146124
rect 252336 146112 252342 146124
rect 259638 146112 259644 146124
rect 252336 146084 259644 146112
rect 252336 146072 252342 146084
rect 259638 146072 259644 146084
rect 259696 146072 259702 146124
rect 324314 145664 324320 145716
rect 324372 145704 324378 145716
rect 327166 145704 327172 145716
rect 324372 145676 327172 145704
rect 324372 145664 324378 145676
rect 327166 145664 327172 145676
rect 327224 145664 327230 145716
rect 253474 145528 253480 145580
rect 253532 145568 253538 145580
rect 307110 145568 307116 145580
rect 253532 145540 307116 145568
rect 253532 145528 253538 145540
rect 307110 145528 307116 145540
rect 307168 145528 307174 145580
rect 184198 144984 184204 145036
rect 184256 145024 184262 145036
rect 213914 145024 213920 145036
rect 184256 144996 213920 145024
rect 184256 144984 184262 144996
rect 213914 144984 213920 144996
rect 213972 144984 213978 145036
rect 303062 144984 303068 145036
rect 303120 145024 303126 145036
rect 307478 145024 307484 145036
rect 303120 144996 307484 145024
rect 303120 144984 303126 144996
rect 307478 144984 307484 144996
rect 307536 144984 307542 145036
rect 174630 144916 174636 144968
rect 174688 144956 174694 144968
rect 214006 144956 214012 144968
rect 174688 144928 214012 144956
rect 174688 144916 174694 144928
rect 214006 144916 214012 144928
rect 214064 144916 214070 144968
rect 279602 144916 279608 144968
rect 279660 144956 279666 144968
rect 307662 144956 307668 144968
rect 279660 144928 307668 144956
rect 279660 144916 279666 144928
rect 307662 144916 307668 144928
rect 307720 144916 307726 144968
rect 252370 144848 252376 144900
rect 252428 144888 252434 144900
rect 267826 144888 267832 144900
rect 252428 144860 267832 144888
rect 252428 144848 252434 144860
rect 267826 144848 267832 144860
rect 267884 144848 267890 144900
rect 324406 144848 324412 144900
rect 324464 144888 324470 144900
rect 338206 144888 338212 144900
rect 324464 144860 338212 144888
rect 324464 144848 324470 144860
rect 338206 144848 338212 144860
rect 338264 144848 338270 144900
rect 252462 144780 252468 144832
rect 252520 144820 252526 144832
rect 262490 144820 262496 144832
rect 252520 144792 262496 144820
rect 252520 144780 252526 144792
rect 262490 144780 262496 144792
rect 262548 144780 262554 144832
rect 324314 144780 324320 144832
rect 324372 144820 324378 144832
rect 336734 144820 336740 144832
rect 324372 144792 336740 144820
rect 324372 144780 324378 144792
rect 336734 144780 336740 144792
rect 336792 144780 336798 144832
rect 290734 144236 290740 144288
rect 290792 144276 290798 144288
rect 307570 144276 307576 144288
rect 290792 144248 307576 144276
rect 290792 144236 290798 144248
rect 307570 144236 307576 144248
rect 307628 144236 307634 144288
rect 253382 144168 253388 144220
rect 253440 144208 253446 144220
rect 307386 144208 307392 144220
rect 253440 144180 307392 144208
rect 253440 144168 253446 144180
rect 307386 144168 307392 144180
rect 307444 144168 307450 144220
rect 304534 143624 304540 143676
rect 304592 143664 304598 143676
rect 307662 143664 307668 143676
rect 304592 143636 307668 143664
rect 304592 143624 304598 143636
rect 307662 143624 307668 143636
rect 307720 143624 307726 143676
rect 167730 143556 167736 143608
rect 167788 143596 167794 143608
rect 213914 143596 213920 143608
rect 167788 143568 213920 143596
rect 167788 143556 167794 143568
rect 213914 143556 213920 143568
rect 213972 143556 213978 143608
rect 257430 143556 257436 143608
rect 257488 143596 257494 143608
rect 306558 143596 306564 143608
rect 257488 143568 306564 143596
rect 257488 143556 257494 143568
rect 306558 143556 306564 143568
rect 306616 143556 306622 143608
rect 252370 143488 252376 143540
rect 252428 143528 252434 143540
rect 264974 143528 264980 143540
rect 252428 143500 264980 143528
rect 252428 143488 252434 143500
rect 264974 143488 264980 143500
rect 265032 143488 265038 143540
rect 324406 143488 324412 143540
rect 324464 143528 324470 143540
rect 345014 143528 345020 143540
rect 324464 143500 345020 143528
rect 324464 143488 324470 143500
rect 345014 143488 345020 143500
rect 345072 143488 345078 143540
rect 252462 143420 252468 143472
rect 252520 143460 252526 143472
rect 263686 143460 263692 143472
rect 252520 143432 263692 143460
rect 252520 143420 252526 143432
rect 263686 143420 263692 143432
rect 263744 143420 263750 143472
rect 324314 143420 324320 143472
rect 324372 143460 324378 143472
rect 343818 143460 343824 143472
rect 324372 143432 343824 143460
rect 324372 143420 324378 143432
rect 343818 143420 343824 143432
rect 343876 143420 343882 143472
rect 251634 143352 251640 143404
rect 251692 143392 251698 143404
rect 255314 143392 255320 143404
rect 251692 143364 255320 143392
rect 251692 143352 251698 143364
rect 255314 143352 255320 143364
rect 255372 143352 255378 143404
rect 322198 142332 322204 142384
rect 322256 142372 322262 142384
rect 324406 142372 324412 142384
rect 322256 142344 324412 142372
rect 322256 142332 322262 142344
rect 324406 142332 324412 142344
rect 324464 142332 324470 142384
rect 202230 142196 202236 142248
rect 202288 142236 202294 142248
rect 213914 142236 213920 142248
rect 202288 142208 213920 142236
rect 202288 142196 202294 142208
rect 213914 142196 213920 142208
rect 213972 142196 213978 142248
rect 276750 142196 276756 142248
rect 276808 142236 276814 142248
rect 307662 142236 307668 142248
rect 276808 142208 307668 142236
rect 276808 142196 276814 142208
rect 307662 142196 307668 142208
rect 307720 142196 307726 142248
rect 173250 142128 173256 142180
rect 173308 142168 173314 142180
rect 214006 142168 214012 142180
rect 173308 142140 214012 142168
rect 173308 142128 173314 142140
rect 214006 142128 214012 142140
rect 214064 142128 214070 142180
rect 253290 142128 253296 142180
rect 253348 142168 253354 142180
rect 307570 142168 307576 142180
rect 253348 142140 307576 142168
rect 253348 142128 253354 142140
rect 307570 142128 307576 142140
rect 307628 142128 307634 142180
rect 324958 142128 324964 142180
rect 325016 142168 325022 142180
rect 325694 142168 325700 142180
rect 325016 142140 325700 142168
rect 325016 142128 325022 142140
rect 325694 142128 325700 142140
rect 325752 142128 325758 142180
rect 252370 142060 252376 142112
rect 252428 142100 252434 142112
rect 271966 142100 271972 142112
rect 252428 142072 271972 142100
rect 252428 142060 252434 142072
rect 271966 142060 271972 142072
rect 272024 142060 272030 142112
rect 324498 142060 324504 142112
rect 324556 142100 324562 142112
rect 352006 142100 352012 142112
rect 324556 142072 352012 142100
rect 324556 142060 324562 142072
rect 352006 142060 352012 142072
rect 352064 142060 352070 142112
rect 324314 141992 324320 142044
rect 324372 142032 324378 142044
rect 346486 142032 346492 142044
rect 324372 142004 346492 142032
rect 324372 141992 324378 142004
rect 346486 141992 346492 142004
rect 346544 141992 346550 142044
rect 294874 141380 294880 141432
rect 294932 141420 294938 141432
rect 306466 141420 306472 141432
rect 294932 141392 306472 141420
rect 294932 141380 294938 141392
rect 306466 141380 306472 141392
rect 306524 141380 306530 141432
rect 252462 141108 252468 141160
rect 252520 141148 252526 141160
rect 259546 141148 259552 141160
rect 252520 141120 259552 141148
rect 252520 141108 252526 141120
rect 259546 141108 259552 141120
rect 259604 141108 259610 141160
rect 210510 140836 210516 140888
rect 210568 140876 210574 140888
rect 214006 140876 214012 140888
rect 210568 140848 214012 140876
rect 210568 140836 210574 140848
rect 214006 140836 214012 140848
rect 214064 140836 214070 140888
rect 171778 140768 171784 140820
rect 171836 140808 171842 140820
rect 213914 140808 213920 140820
rect 171836 140780 213920 140808
rect 171836 140768 171842 140780
rect 213914 140768 213920 140780
rect 213972 140768 213978 140820
rect 251910 140768 251916 140820
rect 251968 140808 251974 140820
rect 254854 140808 254860 140820
rect 251968 140780 254860 140808
rect 251968 140768 251974 140780
rect 254854 140768 254860 140780
rect 254912 140768 254918 140820
rect 252462 140700 252468 140752
rect 252520 140740 252526 140752
rect 281718 140740 281724 140752
rect 252520 140712 281724 140740
rect 252520 140700 252526 140712
rect 281718 140700 281724 140712
rect 281776 140700 281782 140752
rect 324314 140700 324320 140752
rect 324372 140740 324378 140752
rect 328730 140740 328736 140752
rect 324372 140712 328736 140740
rect 324372 140700 324378 140712
rect 328730 140700 328736 140712
rect 328788 140700 328794 140752
rect 252370 140632 252376 140684
rect 252428 140672 252434 140684
rect 256970 140672 256976 140684
rect 252428 140644 256976 140672
rect 252428 140632 252434 140644
rect 256970 140632 256976 140644
rect 257028 140632 257034 140684
rect 180334 140020 180340 140072
rect 180392 140060 180398 140072
rect 214558 140060 214564 140072
rect 180392 140032 214564 140060
rect 180392 140020 180398 140032
rect 214558 140020 214564 140032
rect 214616 140020 214622 140072
rect 252094 140020 252100 140072
rect 252152 140060 252158 140072
rect 290458 140060 290464 140072
rect 252152 140032 290464 140060
rect 252152 140020 252158 140032
rect 290458 140020 290464 140032
rect 290516 140020 290522 140072
rect 282270 139476 282276 139528
rect 282328 139516 282334 139528
rect 307294 139516 307300 139528
rect 282328 139488 307300 139516
rect 282328 139476 282334 139488
rect 307294 139476 307300 139488
rect 307352 139476 307358 139528
rect 207658 139408 207664 139460
rect 207716 139448 207722 139460
rect 213914 139448 213920 139460
rect 207716 139420 213920 139448
rect 207716 139408 207722 139420
rect 213914 139408 213920 139420
rect 213972 139408 213978 139460
rect 267182 139408 267188 139460
rect 267240 139448 267246 139460
rect 307662 139448 307668 139460
rect 267240 139420 307668 139448
rect 267240 139408 267246 139420
rect 307662 139408 307668 139420
rect 307720 139408 307726 139460
rect 252370 139340 252376 139392
rect 252428 139380 252434 139392
rect 274726 139380 274732 139392
rect 252428 139352 274732 139380
rect 252428 139340 252434 139352
rect 274726 139340 274732 139352
rect 274784 139340 274790 139392
rect 324314 139340 324320 139392
rect 324372 139380 324378 139392
rect 343726 139380 343732 139392
rect 324372 139352 343732 139380
rect 324372 139340 324378 139352
rect 343726 139340 343732 139352
rect 343784 139340 343790 139392
rect 252462 139272 252468 139324
rect 252520 139312 252526 139324
rect 262306 139312 262312 139324
rect 252520 139284 262312 139312
rect 252520 139272 252526 139284
rect 262306 139272 262312 139284
rect 262364 139272 262370 139324
rect 324498 139272 324504 139324
rect 324556 139312 324562 139324
rect 341058 139312 341064 139324
rect 324556 139284 341064 139312
rect 324556 139272 324562 139284
rect 341058 139272 341064 139284
rect 341116 139272 341122 139324
rect 294598 138116 294604 138168
rect 294656 138156 294662 138168
rect 307294 138156 307300 138168
rect 294656 138128 307300 138156
rect 294656 138116 294662 138128
rect 307294 138116 307300 138128
rect 307352 138116 307358 138168
rect 278130 138048 278136 138100
rect 278188 138088 278194 138100
rect 307662 138088 307668 138100
rect 278188 138060 307668 138088
rect 278188 138048 278194 138060
rect 307662 138048 307668 138060
rect 307720 138048 307726 138100
rect 196710 137980 196716 138032
rect 196768 138020 196774 138032
rect 213914 138020 213920 138032
rect 196768 137992 213920 138020
rect 196768 137980 196774 137992
rect 213914 137980 213920 137992
rect 213972 137980 213978 138032
rect 250438 137980 250444 138032
rect 250496 138020 250502 138032
rect 307570 138020 307576 138032
rect 250496 137992 307576 138020
rect 250496 137980 250502 137992
rect 307570 137980 307576 137992
rect 307628 137980 307634 138032
rect 252462 137912 252468 137964
rect 252520 137952 252526 137964
rect 276106 137952 276112 137964
rect 252520 137924 276112 137952
rect 252520 137912 252526 137924
rect 276106 137912 276112 137924
rect 276164 137912 276170 137964
rect 324498 137912 324504 137964
rect 324556 137952 324562 137964
rect 335630 137952 335636 137964
rect 324556 137924 335636 137952
rect 324556 137912 324562 137924
rect 335630 137912 335636 137924
rect 335688 137912 335694 137964
rect 252370 137844 252376 137896
rect 252428 137884 252434 137896
rect 273438 137884 273444 137896
rect 252428 137856 273444 137884
rect 252428 137844 252434 137856
rect 273438 137844 273444 137856
rect 273496 137844 273502 137896
rect 324314 137844 324320 137896
rect 324372 137884 324378 137896
rect 334158 137884 334164 137896
rect 324372 137856 334164 137884
rect 324372 137844 324378 137856
rect 334158 137844 334164 137856
rect 334216 137844 334222 137896
rect 177574 137232 177580 137284
rect 177632 137272 177638 137284
rect 214558 137272 214564 137284
rect 177632 137244 214564 137272
rect 177632 137232 177638 137244
rect 214558 137232 214564 137244
rect 214616 137232 214622 137284
rect 254854 137232 254860 137284
rect 254912 137272 254918 137284
rect 307018 137272 307024 137284
rect 254912 137244 307024 137272
rect 254912 137232 254918 137244
rect 307018 137232 307024 137244
rect 307076 137232 307082 137284
rect 2774 136960 2780 137012
rect 2832 137000 2838 137012
rect 4798 137000 4804 137012
rect 2832 136972 4804 137000
rect 2832 136960 2838 136972
rect 4798 136960 4804 136972
rect 4856 136960 4862 137012
rect 292022 136688 292028 136740
rect 292080 136728 292086 136740
rect 307570 136728 307576 136740
rect 292080 136700 307576 136728
rect 292080 136688 292086 136700
rect 307570 136688 307576 136700
rect 307628 136688 307634 136740
rect 166258 136620 166264 136672
rect 166316 136660 166322 136672
rect 213914 136660 213920 136672
rect 166316 136632 213920 136660
rect 166316 136620 166322 136632
rect 213914 136620 213920 136632
rect 213972 136620 213978 136672
rect 250530 136620 250536 136672
rect 250588 136660 250594 136672
rect 307662 136660 307668 136672
rect 250588 136632 307668 136660
rect 250588 136620 250594 136632
rect 307662 136620 307668 136632
rect 307720 136620 307726 136672
rect 252278 136552 252284 136604
rect 252336 136592 252342 136604
rect 291930 136592 291936 136604
rect 252336 136564 291936 136592
rect 252336 136552 252342 136564
rect 291930 136552 291936 136564
rect 291988 136552 291994 136604
rect 324498 136552 324504 136604
rect 324556 136592 324562 136604
rect 342254 136592 342260 136604
rect 324556 136564 342260 136592
rect 324556 136552 324562 136564
rect 342254 136552 342260 136564
rect 342312 136552 342318 136604
rect 252462 136484 252468 136536
rect 252520 136524 252526 136536
rect 289170 136524 289176 136536
rect 252520 136496 289176 136524
rect 252520 136484 252526 136496
rect 289170 136484 289176 136496
rect 289228 136484 289234 136536
rect 252370 136416 252376 136468
rect 252428 136456 252434 136468
rect 269758 136456 269764 136468
rect 252428 136428 269764 136456
rect 252428 136416 252434 136428
rect 269758 136416 269764 136428
rect 269816 136416 269822 136468
rect 252002 136348 252008 136400
rect 252060 136388 252066 136400
rect 254578 136388 254584 136400
rect 252060 136360 254584 136388
rect 252060 136348 252066 136360
rect 254578 136348 254584 136360
rect 254636 136348 254642 136400
rect 324314 136348 324320 136400
rect 324372 136388 324378 136400
rect 327258 136388 327264 136400
rect 324372 136360 327264 136388
rect 324372 136348 324378 136360
rect 327258 136348 327264 136360
rect 327316 136348 327322 136400
rect 300210 135464 300216 135516
rect 300268 135504 300274 135516
rect 306742 135504 306748 135516
rect 300268 135476 306748 135504
rect 300268 135464 300274 135476
rect 306742 135464 306748 135476
rect 306800 135464 306806 135516
rect 289262 135396 289268 135448
rect 289320 135436 289326 135448
rect 307662 135436 307668 135448
rect 289320 135408 307668 135436
rect 289320 135396 289326 135408
rect 307662 135396 307668 135408
rect 307720 135396 307726 135448
rect 285030 135328 285036 135380
rect 285088 135368 285094 135380
rect 307478 135368 307484 135380
rect 285088 135340 307484 135368
rect 285088 135328 285094 135340
rect 307478 135328 307484 135340
rect 307536 135328 307542 135380
rect 178770 135260 178776 135312
rect 178828 135300 178834 135312
rect 213914 135300 213920 135312
rect 178828 135272 213920 135300
rect 178828 135260 178834 135272
rect 213914 135260 213920 135272
rect 213972 135260 213978 135312
rect 265710 135260 265716 135312
rect 265768 135300 265774 135312
rect 307570 135300 307576 135312
rect 265768 135272 307576 135300
rect 265768 135260 265774 135272
rect 307570 135260 307576 135272
rect 307628 135260 307634 135312
rect 252370 135192 252376 135244
rect 252428 135232 252434 135244
rect 295978 135232 295984 135244
rect 252428 135204 295984 135232
rect 252428 135192 252434 135204
rect 295978 135192 295984 135204
rect 296036 135192 296042 135244
rect 324314 135192 324320 135244
rect 324372 135232 324378 135244
rect 331398 135232 331404 135244
rect 324372 135204 331404 135232
rect 324372 135192 324378 135204
rect 331398 135192 331404 135204
rect 331456 135192 331462 135244
rect 252462 135124 252468 135176
rect 252520 135164 252526 135176
rect 289078 135164 289084 135176
rect 252520 135136 289084 135164
rect 252520 135124 252526 135136
rect 289078 135124 289084 135136
rect 289136 135124 289142 135176
rect 286686 134512 286692 134564
rect 286744 134552 286750 134564
rect 307386 134552 307392 134564
rect 286744 134524 307392 134552
rect 286744 134512 286750 134524
rect 307386 134512 307392 134524
rect 307444 134512 307450 134564
rect 181438 133900 181444 133952
rect 181496 133940 181502 133952
rect 213914 133940 213920 133952
rect 181496 133912 213920 133940
rect 181496 133900 181502 133912
rect 213914 133900 213920 133912
rect 213972 133900 213978 133952
rect 293218 133900 293224 133952
rect 293276 133940 293282 133952
rect 307662 133940 307668 133952
rect 293276 133912 307668 133940
rect 293276 133900 293282 133912
rect 307662 133900 307668 133912
rect 307720 133900 307726 133952
rect 252370 133832 252376 133884
rect 252428 133872 252434 133884
rect 296070 133872 296076 133884
rect 252428 133844 296076 133872
rect 252428 133832 252434 133844
rect 296070 133832 296076 133844
rect 296128 133832 296134 133884
rect 324314 133832 324320 133884
rect 324372 133872 324378 133884
rect 345198 133872 345204 133884
rect 324372 133844 345204 133872
rect 324372 133832 324378 133844
rect 345198 133832 345204 133844
rect 345256 133832 345262 133884
rect 252278 133764 252284 133816
rect 252336 133804 252342 133816
rect 268378 133804 268384 133816
rect 252336 133776 268384 133804
rect 252336 133764 252342 133776
rect 268378 133764 268384 133776
rect 268436 133764 268442 133816
rect 252462 133696 252468 133748
rect 252520 133736 252526 133748
rect 266998 133736 267004 133748
rect 252520 133708 267004 133736
rect 252520 133696 252526 133708
rect 266998 133696 267004 133708
rect 267056 133696 267062 133748
rect 295978 132608 295984 132660
rect 296036 132648 296042 132660
rect 306558 132648 306564 132660
rect 296036 132620 306564 132648
rect 296036 132608 296042 132620
rect 306558 132608 306564 132620
rect 306616 132608 306622 132660
rect 202322 132540 202328 132592
rect 202380 132580 202386 132592
rect 214006 132580 214012 132592
rect 202380 132552 214012 132580
rect 202380 132540 202386 132552
rect 214006 132540 214012 132552
rect 214064 132540 214070 132592
rect 287790 132540 287796 132592
rect 287848 132580 287854 132592
rect 307110 132580 307116 132592
rect 287848 132552 307116 132580
rect 287848 132540 287854 132552
rect 307110 132540 307116 132552
rect 307168 132540 307174 132592
rect 173342 132472 173348 132524
rect 173400 132512 173406 132524
rect 213914 132512 213920 132524
rect 173400 132484 213920 132512
rect 173400 132472 173406 132484
rect 213914 132472 213920 132484
rect 213972 132472 213978 132524
rect 273898 132472 273904 132524
rect 273956 132512 273962 132524
rect 307662 132512 307668 132524
rect 273956 132484 307668 132512
rect 273956 132472 273962 132484
rect 307662 132472 307668 132484
rect 307720 132472 307726 132524
rect 252278 132404 252284 132456
rect 252336 132444 252342 132456
rect 300118 132444 300124 132456
rect 252336 132416 300124 132444
rect 252336 132404 252342 132416
rect 300118 132404 300124 132416
rect 300176 132404 300182 132456
rect 252370 132336 252376 132388
rect 252428 132376 252434 132388
rect 286410 132376 286416 132388
rect 252428 132348 286416 132376
rect 252428 132336 252434 132348
rect 286410 132336 286416 132348
rect 286468 132336 286474 132388
rect 252462 132268 252468 132320
rect 252520 132308 252526 132320
rect 264422 132308 264428 132320
rect 252520 132280 264428 132308
rect 252520 132268 252526 132280
rect 264422 132268 264428 132280
rect 264480 132268 264486 132320
rect 203610 131180 203616 131232
rect 203668 131220 203674 131232
rect 214006 131220 214012 131232
rect 203668 131192 214012 131220
rect 203668 131180 203674 131192
rect 214006 131180 214012 131192
rect 214064 131180 214070 131232
rect 286502 131180 286508 131232
rect 286560 131220 286566 131232
rect 306926 131220 306932 131232
rect 286560 131192 306932 131220
rect 286560 131180 286566 131192
rect 306926 131180 306932 131192
rect 306984 131180 306990 131232
rect 171870 131112 171876 131164
rect 171928 131152 171934 131164
rect 213914 131152 213920 131164
rect 171928 131124 213920 131152
rect 171928 131112 171934 131124
rect 213914 131112 213920 131124
rect 213972 131112 213978 131164
rect 283558 131112 283564 131164
rect 283616 131152 283622 131164
rect 306558 131152 306564 131164
rect 283616 131124 306564 131152
rect 283616 131112 283622 131124
rect 306558 131112 306564 131124
rect 306616 131112 306622 131164
rect 252462 131044 252468 131096
rect 252520 131084 252526 131096
rect 275370 131084 275376 131096
rect 252520 131056 275376 131084
rect 252520 131044 252526 131056
rect 275370 131044 275376 131056
rect 275428 131044 275434 131096
rect 324314 131044 324320 131096
rect 324372 131084 324378 131096
rect 347866 131084 347872 131096
rect 324372 131056 347872 131084
rect 324372 131044 324378 131056
rect 347866 131044 347872 131056
rect 347924 131044 347930 131096
rect 252370 130976 252376 131028
rect 252428 131016 252434 131028
rect 269850 131016 269856 131028
rect 252428 130988 269856 131016
rect 252428 130976 252434 130988
rect 269850 130976 269856 130988
rect 269908 130976 269914 131028
rect 324406 130976 324412 131028
rect 324464 131016 324470 131028
rect 330018 131016 330024 131028
rect 324464 130988 330024 131016
rect 324464 130976 324470 130988
rect 330018 130976 330024 130988
rect 330076 130976 330082 131028
rect 252278 130908 252284 130960
rect 252336 130948 252342 130960
rect 262858 130948 262864 130960
rect 252336 130920 262864 130948
rect 252336 130908 252342 130920
rect 262858 130908 262864 130920
rect 262916 130908 262922 130960
rect 269942 130364 269948 130416
rect 270000 130404 270006 130416
rect 307294 130404 307300 130416
rect 270000 130376 307300 130404
rect 270000 130364 270006 130376
rect 307294 130364 307300 130376
rect 307352 130364 307358 130416
rect 290642 129820 290648 129872
rect 290700 129860 290706 129872
rect 307478 129860 307484 129872
rect 290700 129832 307484 129860
rect 290700 129820 290706 129832
rect 307478 129820 307484 129832
rect 307536 129820 307542 129872
rect 171962 129752 171968 129804
rect 172020 129792 172026 129804
rect 213914 129792 213920 129804
rect 172020 129764 213920 129792
rect 172020 129752 172026 129764
rect 213914 129752 213920 129764
rect 213972 129752 213978 129804
rect 275278 129752 275284 129804
rect 275336 129792 275342 129804
rect 307662 129792 307668 129804
rect 275336 129764 307668 129792
rect 275336 129752 275342 129764
rect 307662 129752 307668 129764
rect 307720 129752 307726 129804
rect 252370 129684 252376 129736
rect 252428 129724 252434 129736
rect 276658 129724 276664 129736
rect 252428 129696 276664 129724
rect 252428 129684 252434 129696
rect 276658 129684 276664 129696
rect 276716 129684 276722 129736
rect 324314 129684 324320 129736
rect 324372 129724 324378 129736
rect 329926 129724 329932 129736
rect 324372 129696 329932 129724
rect 324372 129684 324378 129696
rect 329926 129684 329932 129696
rect 329984 129684 329990 129736
rect 252462 129616 252468 129668
rect 252520 129656 252526 129668
rect 271322 129656 271328 129668
rect 252520 129628 271328 129656
rect 252520 129616 252526 129628
rect 271322 129616 271328 129628
rect 271380 129616 271386 129668
rect 324406 129616 324412 129668
rect 324464 129656 324470 129668
rect 329834 129656 329840 129668
rect 324464 129628 329840 129656
rect 324464 129616 324470 129628
rect 329834 129616 329840 129628
rect 329892 129616 329898 129668
rect 290550 128460 290556 128512
rect 290608 128500 290614 128512
rect 307478 128500 307484 128512
rect 290608 128472 307484 128500
rect 290608 128460 290614 128472
rect 307478 128460 307484 128472
rect 307536 128460 307542 128512
rect 280890 128392 280896 128444
rect 280948 128432 280954 128444
rect 307570 128432 307576 128444
rect 280948 128404 307576 128432
rect 280948 128392 280954 128404
rect 307570 128392 307576 128404
rect 307628 128392 307634 128444
rect 176010 128324 176016 128376
rect 176068 128364 176074 128376
rect 213914 128364 213920 128376
rect 176068 128336 213920 128364
rect 176068 128324 176074 128336
rect 213914 128324 213920 128336
rect 213972 128324 213978 128376
rect 252186 128324 252192 128376
rect 252244 128364 252250 128376
rect 260190 128364 260196 128376
rect 252244 128336 260196 128364
rect 252244 128324 252250 128336
rect 260190 128324 260196 128336
rect 260248 128324 260254 128376
rect 271138 128324 271144 128376
rect 271196 128364 271202 128376
rect 307662 128364 307668 128376
rect 271196 128336 307668 128364
rect 271196 128324 271202 128336
rect 307662 128324 307668 128336
rect 307720 128324 307726 128376
rect 252462 128256 252468 128308
rect 252520 128296 252526 128308
rect 283742 128296 283748 128308
rect 252520 128268 283748 128296
rect 252520 128256 252526 128268
rect 283742 128256 283748 128268
rect 283800 128256 283806 128308
rect 324314 128256 324320 128308
rect 324372 128296 324378 128308
rect 328546 128296 328552 128308
rect 324372 128268 328552 128296
rect 324372 128256 324378 128268
rect 328546 128256 328552 128268
rect 328604 128256 328610 128308
rect 252278 128188 252284 128240
rect 252336 128228 252342 128240
rect 281074 128228 281080 128240
rect 252336 128200 281080 128228
rect 252336 128188 252342 128200
rect 281074 128188 281080 128200
rect 281132 128188 281138 128240
rect 252370 128120 252376 128172
rect 252428 128160 252434 128172
rect 278222 128160 278228 128172
rect 252428 128132 278228 128160
rect 252428 128120 252434 128132
rect 278222 128120 278228 128132
rect 278280 128120 278286 128172
rect 283650 127100 283656 127152
rect 283708 127140 283714 127152
rect 307570 127140 307576 127152
rect 283708 127112 307576 127140
rect 283708 127100 283714 127112
rect 307570 127100 307576 127112
rect 307628 127100 307634 127152
rect 282178 127032 282184 127084
rect 282236 127072 282242 127084
rect 307662 127072 307668 127084
rect 282236 127044 307668 127072
rect 282236 127032 282242 127044
rect 307662 127032 307668 127044
rect 307720 127032 307726 127084
rect 198090 126964 198096 127016
rect 198148 127004 198154 127016
rect 213914 127004 213920 127016
rect 198148 126976 213920 127004
rect 198148 126964 198154 126976
rect 213914 126964 213920 126976
rect 213972 126964 213978 127016
rect 280982 126964 280988 127016
rect 281040 127004 281046 127016
rect 307478 127004 307484 127016
rect 281040 126976 307484 127004
rect 281040 126964 281046 126976
rect 307478 126964 307484 126976
rect 307536 126964 307542 127016
rect 252462 126896 252468 126948
rect 252520 126936 252526 126948
rect 302878 126936 302884 126948
rect 252520 126908 302884 126936
rect 252520 126896 252526 126908
rect 302878 126896 302884 126908
rect 302936 126896 302942 126948
rect 251726 126828 251732 126880
rect 251784 126868 251790 126880
rect 254854 126868 254860 126880
rect 251784 126840 254860 126868
rect 251784 126828 251790 126840
rect 254854 126828 254860 126840
rect 254912 126828 254918 126880
rect 252278 126216 252284 126268
rect 252336 126256 252342 126268
rect 305730 126256 305736 126268
rect 252336 126228 305736 126256
rect 252336 126216 252342 126228
rect 305730 126216 305736 126228
rect 305788 126216 305794 126268
rect 207750 125672 207756 125724
rect 207808 125712 207814 125724
rect 213914 125712 213920 125724
rect 207808 125684 213920 125712
rect 207808 125672 207814 125684
rect 213914 125672 213920 125684
rect 213972 125672 213978 125724
rect 289354 125672 289360 125724
rect 289412 125712 289418 125724
rect 306558 125712 306564 125724
rect 289412 125684 306564 125712
rect 289412 125672 289418 125684
rect 306558 125672 306564 125684
rect 306616 125672 306622 125724
rect 59262 125604 59268 125656
rect 59320 125644 59326 125656
rect 65150 125644 65156 125656
rect 59320 125616 65156 125644
rect 59320 125604 59326 125616
rect 65150 125604 65156 125616
rect 65208 125604 65214 125656
rect 176102 125604 176108 125656
rect 176160 125644 176166 125656
rect 214006 125644 214012 125656
rect 176160 125616 214012 125644
rect 176160 125604 176166 125616
rect 214006 125604 214012 125616
rect 214064 125604 214070 125656
rect 254578 125604 254584 125656
rect 254636 125644 254642 125656
rect 307662 125644 307668 125656
rect 254636 125616 307668 125644
rect 254636 125604 254642 125616
rect 307662 125604 307668 125616
rect 307720 125604 307726 125656
rect 252462 125536 252468 125588
rect 252520 125576 252526 125588
rect 298830 125576 298836 125588
rect 252520 125548 298836 125576
rect 252520 125536 252526 125548
rect 298830 125536 298836 125548
rect 298888 125536 298894 125588
rect 324314 125536 324320 125588
rect 324372 125576 324378 125588
rect 332686 125576 332692 125588
rect 324372 125548 332692 125576
rect 324372 125536 324378 125548
rect 332686 125536 332692 125548
rect 332744 125536 332750 125588
rect 252370 125468 252376 125520
rect 252428 125508 252434 125520
rect 287974 125508 287980 125520
rect 252428 125480 287980 125508
rect 252428 125468 252434 125480
rect 287974 125468 287980 125480
rect 288032 125468 288038 125520
rect 302878 124380 302884 124432
rect 302936 124420 302942 124432
rect 307662 124420 307668 124432
rect 302936 124392 307668 124420
rect 302936 124380 302942 124392
rect 307662 124380 307668 124392
rect 307720 124380 307726 124432
rect 298738 124312 298744 124364
rect 298796 124352 298802 124364
rect 306558 124352 306564 124364
rect 298796 124324 306564 124352
rect 298796 124312 298802 124324
rect 306558 124312 306564 124324
rect 306616 124312 306622 124364
rect 187142 124244 187148 124296
rect 187200 124284 187206 124296
rect 213914 124284 213920 124296
rect 187200 124256 213920 124284
rect 187200 124244 187206 124256
rect 213914 124244 213920 124256
rect 213972 124244 213978 124296
rect 287882 124244 287888 124296
rect 287940 124284 287946 124296
rect 307478 124284 307484 124296
rect 287940 124256 307484 124284
rect 287940 124244 287946 124256
rect 307478 124244 307484 124256
rect 307536 124244 307542 124296
rect 62022 124176 62028 124228
rect 62080 124216 62086 124228
rect 65518 124216 65524 124228
rect 62080 124188 65524 124216
rect 62080 124176 62086 124188
rect 65518 124176 65524 124188
rect 65576 124176 65582 124228
rect 169202 124176 169208 124228
rect 169260 124216 169266 124228
rect 214006 124216 214012 124228
rect 169260 124188 214012 124216
rect 169260 124176 169266 124188
rect 214006 124176 214012 124188
rect 214064 124176 214070 124228
rect 255958 124176 255964 124228
rect 256016 124216 256022 124228
rect 307570 124216 307576 124228
rect 256016 124188 307576 124216
rect 256016 124176 256022 124188
rect 307570 124176 307576 124188
rect 307628 124176 307634 124228
rect 252462 124108 252468 124160
rect 252520 124148 252526 124160
rect 301498 124148 301504 124160
rect 252520 124120 301504 124148
rect 252520 124108 252526 124120
rect 301498 124108 301504 124120
rect 301556 124108 301562 124160
rect 324314 124108 324320 124160
rect 324372 124148 324378 124160
rect 340966 124148 340972 124160
rect 324372 124120 340972 124148
rect 324372 124108 324378 124120
rect 340966 124108 340972 124120
rect 341024 124108 341030 124160
rect 252370 124040 252376 124092
rect 252428 124080 252434 124092
rect 271230 124080 271236 124092
rect 252428 124052 271236 124080
rect 252428 124040 252434 124052
rect 271230 124040 271236 124052
rect 271288 124040 271294 124092
rect 324406 124040 324412 124092
rect 324464 124080 324470 124092
rect 338390 124080 338396 124092
rect 324464 124052 338396 124080
rect 324464 124040 324470 124052
rect 338390 124040 338396 124052
rect 338448 124040 338454 124092
rect 252278 123972 252284 124024
rect 252336 124012 252342 124024
rect 257522 124012 257528 124024
rect 252336 123984 257528 124012
rect 252336 123972 252342 123984
rect 257522 123972 257528 123984
rect 257580 123972 257586 124024
rect 301682 122952 301688 123004
rect 301740 122992 301746 123004
rect 307662 122992 307668 123004
rect 301740 122964 307668 122992
rect 301740 122952 301746 122964
rect 307662 122952 307668 122964
rect 307720 122952 307726 123004
rect 170582 122884 170588 122936
rect 170640 122924 170646 122936
rect 213914 122924 213920 122936
rect 170640 122896 213920 122924
rect 170640 122884 170646 122896
rect 213914 122884 213920 122896
rect 213972 122884 213978 122936
rect 289078 122884 289084 122936
rect 289136 122924 289142 122936
rect 307478 122924 307484 122936
rect 289136 122896 307484 122924
rect 289136 122884 289142 122896
rect 307478 122884 307484 122896
rect 307536 122884 307542 122936
rect 61930 122816 61936 122868
rect 61988 122856 61994 122868
rect 66070 122856 66076 122868
rect 61988 122828 66076 122856
rect 61988 122816 61994 122828
rect 66070 122816 66076 122828
rect 66128 122816 66134 122868
rect 169110 122816 169116 122868
rect 169168 122856 169174 122868
rect 214006 122856 214012 122868
rect 169168 122828 214012 122856
rect 169168 122816 169174 122828
rect 214006 122816 214012 122828
rect 214064 122816 214070 122868
rect 272518 122816 272524 122868
rect 272576 122856 272582 122868
rect 307570 122856 307576 122868
rect 272576 122828 307576 122856
rect 272576 122816 272582 122828
rect 307570 122816 307576 122828
rect 307628 122816 307634 122868
rect 252462 122748 252468 122800
rect 252520 122788 252526 122800
rect 297450 122788 297456 122800
rect 252520 122760 297456 122788
rect 252520 122748 252526 122760
rect 297450 122748 297456 122760
rect 297508 122748 297514 122800
rect 324314 122748 324320 122800
rect 324372 122788 324378 122800
rect 358814 122788 358820 122800
rect 324372 122760 358820 122788
rect 324372 122748 324378 122760
rect 358814 122748 358820 122760
rect 358872 122748 358878 122800
rect 252278 122680 252284 122732
rect 252336 122720 252342 122732
rect 264238 122720 264244 122732
rect 252336 122692 264244 122720
rect 252336 122680 252342 122692
rect 264238 122680 264244 122692
rect 264296 122680 264302 122732
rect 252370 122408 252376 122460
rect 252428 122448 252434 122460
rect 258902 122448 258908 122460
rect 252428 122420 258908 122448
rect 252428 122408 252434 122420
rect 258902 122408 258908 122420
rect 258960 122408 258966 122460
rect 297358 121592 297364 121644
rect 297416 121632 297422 121644
rect 307478 121632 307484 121644
rect 297416 121604 307484 121632
rect 297416 121592 297422 121604
rect 307478 121592 307484 121604
rect 307536 121592 307542 121644
rect 209222 121524 209228 121576
rect 209280 121564 209286 121576
rect 214006 121564 214012 121576
rect 209280 121536 214012 121564
rect 209280 121524 209286 121536
rect 214006 121524 214012 121536
rect 214064 121524 214070 121576
rect 293310 121524 293316 121576
rect 293368 121564 293374 121576
rect 307570 121564 307576 121576
rect 293368 121536 307576 121564
rect 293368 121524 293374 121536
rect 307570 121524 307576 121536
rect 307628 121524 307634 121576
rect 177390 121456 177396 121508
rect 177448 121496 177454 121508
rect 213914 121496 213920 121508
rect 177448 121468 213920 121496
rect 177448 121456 177454 121468
rect 213914 121456 213920 121468
rect 213972 121456 213978 121508
rect 266998 121456 267004 121508
rect 267056 121496 267062 121508
rect 307662 121496 307668 121508
rect 267056 121468 307668 121496
rect 267056 121456 267062 121468
rect 307662 121456 307668 121468
rect 307720 121456 307726 121508
rect 252370 121388 252376 121440
rect 252428 121428 252434 121440
rect 291838 121428 291844 121440
rect 252428 121400 291844 121428
rect 252428 121388 252434 121400
rect 291838 121388 291844 121400
rect 291896 121388 291902 121440
rect 324314 121388 324320 121440
rect 324372 121428 324378 121440
rect 356054 121428 356060 121440
rect 324372 121400 356060 121428
rect 324372 121388 324378 121400
rect 356054 121388 356060 121400
rect 356112 121388 356118 121440
rect 252462 121320 252468 121372
rect 252520 121360 252526 121372
rect 265618 121360 265624 121372
rect 252520 121332 265624 121360
rect 252520 121320 252526 121332
rect 265618 121320 265624 121332
rect 265676 121320 265682 121372
rect 252462 120912 252468 120964
rect 252520 120952 252526 120964
rect 258718 120952 258724 120964
rect 252520 120924 258724 120952
rect 252520 120912 252526 120924
rect 258718 120912 258724 120924
rect 258776 120912 258782 120964
rect 296070 120232 296076 120284
rect 296128 120272 296134 120284
rect 307662 120272 307668 120284
rect 296128 120244 307668 120272
rect 296128 120232 296134 120244
rect 307662 120232 307668 120244
rect 307720 120232 307726 120284
rect 188430 120164 188436 120216
rect 188488 120204 188494 120216
rect 213914 120204 213920 120216
rect 188488 120176 213920 120204
rect 188488 120164 188494 120176
rect 213914 120164 213920 120176
rect 213972 120164 213978 120216
rect 286410 120164 286416 120216
rect 286468 120204 286474 120216
rect 307570 120204 307576 120216
rect 286468 120176 307576 120204
rect 286468 120164 286474 120176
rect 307570 120164 307576 120176
rect 307628 120164 307634 120216
rect 166350 120096 166356 120148
rect 166408 120136 166414 120148
rect 214006 120136 214012 120148
rect 166408 120108 214012 120136
rect 166408 120096 166414 120108
rect 214006 120096 214012 120108
rect 214064 120096 214070 120148
rect 271230 120096 271236 120148
rect 271288 120136 271294 120148
rect 307110 120136 307116 120148
rect 271288 120108 307116 120136
rect 271288 120096 271294 120108
rect 307110 120096 307116 120108
rect 307168 120096 307174 120148
rect 252462 120028 252468 120080
rect 252520 120068 252526 120080
rect 262950 120068 262956 120080
rect 252520 120040 262956 120068
rect 252520 120028 252526 120040
rect 262950 120028 262956 120040
rect 263008 120028 263014 120080
rect 252278 119960 252284 120012
rect 252336 120000 252342 120012
rect 253474 120000 253480 120012
rect 252336 119972 253480 120000
rect 252336 119960 252342 119972
rect 253474 119960 253480 119972
rect 253532 119960 253538 120012
rect 252370 119348 252376 119400
rect 252428 119388 252434 119400
rect 293402 119388 293408 119400
rect 252428 119360 293408 119388
rect 252428 119348 252434 119360
rect 293402 119348 293408 119360
rect 293460 119348 293466 119400
rect 170398 118804 170404 118856
rect 170456 118844 170462 118856
rect 213914 118844 213920 118856
rect 170456 118816 213920 118844
rect 170456 118804 170462 118816
rect 213914 118804 213920 118816
rect 213972 118804 213978 118856
rect 304258 118804 304264 118856
rect 304316 118844 304322 118856
rect 307662 118844 307668 118856
rect 304316 118816 307668 118844
rect 304316 118804 304322 118816
rect 307662 118804 307668 118816
rect 307720 118804 307726 118856
rect 185670 118736 185676 118788
rect 185728 118776 185734 118788
rect 214006 118776 214012 118788
rect 185728 118748 214012 118776
rect 185728 118736 185734 118748
rect 214006 118736 214012 118748
rect 214064 118736 214070 118788
rect 291838 118736 291844 118788
rect 291896 118776 291902 118788
rect 307570 118776 307576 118788
rect 291896 118748 307576 118776
rect 291896 118736 291902 118748
rect 307570 118736 307576 118748
rect 307628 118736 307634 118788
rect 262858 118668 262864 118720
rect 262916 118708 262922 118720
rect 307110 118708 307116 118720
rect 262916 118680 307116 118708
rect 262916 118668 262922 118680
rect 307110 118668 307116 118680
rect 307168 118668 307174 118720
rect 252462 118600 252468 118652
rect 252520 118640 252526 118652
rect 264330 118640 264336 118652
rect 252520 118612 264336 118640
rect 252520 118600 252526 118612
rect 264330 118600 264336 118612
rect 264388 118600 264394 118652
rect 324406 118600 324412 118652
rect 324464 118640 324470 118652
rect 345106 118640 345112 118652
rect 324464 118612 345112 118640
rect 324464 118600 324470 118612
rect 345106 118600 345112 118612
rect 345164 118600 345170 118652
rect 324314 118532 324320 118584
rect 324372 118572 324378 118584
rect 339678 118572 339684 118584
rect 324372 118544 339684 118572
rect 324372 118532 324378 118544
rect 339678 118532 339684 118544
rect 339736 118532 339742 118584
rect 252462 117648 252468 117700
rect 252520 117688 252526 117700
rect 258810 117688 258816 117700
rect 252520 117660 258816 117688
rect 252520 117648 252526 117660
rect 258810 117648 258816 117660
rect 258868 117648 258874 117700
rect 300118 117512 300124 117564
rect 300176 117552 300182 117564
rect 306558 117552 306564 117564
rect 300176 117524 306564 117552
rect 300176 117512 300182 117524
rect 306558 117512 306564 117524
rect 306616 117512 306622 117564
rect 298830 117444 298836 117496
rect 298888 117484 298894 117496
rect 307662 117484 307668 117496
rect 298888 117456 307668 117484
rect 298888 117444 298894 117456
rect 307662 117444 307668 117456
rect 307720 117444 307726 117496
rect 174722 117376 174728 117428
rect 174780 117416 174786 117428
rect 214006 117416 214012 117428
rect 174780 117388 214012 117416
rect 174780 117376 174786 117388
rect 214006 117376 214012 117388
rect 214064 117376 214070 117428
rect 265618 117376 265624 117428
rect 265676 117416 265682 117428
rect 307570 117416 307576 117428
rect 265676 117388 307576 117416
rect 265676 117376 265682 117388
rect 307570 117376 307576 117388
rect 307628 117376 307634 117428
rect 170674 117308 170680 117360
rect 170732 117348 170738 117360
rect 213914 117348 213920 117360
rect 170732 117320 213920 117348
rect 170732 117308 170738 117320
rect 213914 117308 213920 117320
rect 213972 117308 213978 117360
rect 264238 117308 264244 117360
rect 264296 117348 264302 117360
rect 307110 117348 307116 117360
rect 264296 117320 307116 117348
rect 264296 117308 264302 117320
rect 307110 117308 307116 117320
rect 307168 117308 307174 117360
rect 252462 117240 252468 117292
rect 252520 117280 252526 117292
rect 282454 117280 282460 117292
rect 252520 117252 282460 117280
rect 252520 117240 252526 117252
rect 282454 117240 282460 117252
rect 282512 117240 282518 117292
rect 324314 117240 324320 117292
rect 324372 117280 324378 117292
rect 338298 117280 338304 117292
rect 324372 117252 338304 117280
rect 324372 117240 324378 117252
rect 338298 117240 338304 117252
rect 338356 117240 338362 117292
rect 252370 117172 252376 117224
rect 252428 117212 252434 117224
rect 268470 117212 268476 117224
rect 252428 117184 268476 117212
rect 252428 117172 252434 117184
rect 268470 117172 268476 117184
rect 268528 117172 268534 117224
rect 296346 116560 296352 116612
rect 296404 116600 296410 116612
rect 307018 116600 307024 116612
rect 296404 116572 307024 116600
rect 296404 116560 296410 116572
rect 307018 116560 307024 116572
rect 307076 116560 307082 116612
rect 252462 116492 252468 116544
rect 252520 116532 252526 116544
rect 260098 116532 260104 116544
rect 252520 116504 260104 116532
rect 252520 116492 252526 116504
rect 260098 116492 260104 116504
rect 260156 116492 260162 116544
rect 198182 116016 198188 116068
rect 198240 116056 198246 116068
rect 214006 116056 214012 116068
rect 198240 116028 214012 116056
rect 198240 116016 198246 116028
rect 214006 116016 214012 116028
rect 214064 116016 214070 116068
rect 282362 116016 282368 116068
rect 282420 116056 282426 116068
rect 306926 116056 306932 116068
rect 282420 116028 306932 116056
rect 282420 116016 282426 116028
rect 306926 116016 306932 116028
rect 306984 116016 306990 116068
rect 181530 115948 181536 116000
rect 181588 115988 181594 116000
rect 213914 115988 213920 116000
rect 181588 115960 213920 115988
rect 181588 115948 181594 115960
rect 213914 115948 213920 115960
rect 213972 115948 213978 116000
rect 268378 115948 268384 116000
rect 268436 115988 268442 116000
rect 307662 115988 307668 116000
rect 268436 115960 307668 115988
rect 268436 115948 268442 115960
rect 307662 115948 307668 115960
rect 307720 115948 307726 116000
rect 252370 115880 252376 115932
rect 252428 115920 252434 115932
rect 267090 115920 267096 115932
rect 252428 115892 267096 115920
rect 252428 115880 252434 115892
rect 267090 115880 267096 115892
rect 267148 115880 267154 115932
rect 324406 115880 324412 115932
rect 324464 115920 324470 115932
rect 351914 115920 351920 115932
rect 324464 115892 351920 115920
rect 324464 115880 324470 115892
rect 351914 115880 351920 115892
rect 351972 115880 351978 115932
rect 324314 115812 324320 115864
rect 324372 115852 324378 115864
rect 342438 115852 342444 115864
rect 324372 115824 342444 115852
rect 324372 115812 324378 115824
rect 342438 115812 342444 115824
rect 342496 115812 342502 115864
rect 169018 115268 169024 115320
rect 169076 115308 169082 115320
rect 203518 115308 203524 115320
rect 169076 115280 203524 115308
rect 169076 115268 169082 115280
rect 203518 115268 203524 115280
rect 203576 115268 203582 115320
rect 173434 115200 173440 115252
rect 173492 115240 173498 115252
rect 214650 115240 214656 115252
rect 173492 115212 214656 115240
rect 173492 115200 173498 115212
rect 214650 115200 214656 115212
rect 214708 115200 214714 115252
rect 252462 115200 252468 115252
rect 252520 115240 252526 115252
rect 297634 115240 297640 115252
rect 252520 115212 297640 115240
rect 252520 115200 252526 115212
rect 297634 115200 297640 115212
rect 297692 115200 297698 115252
rect 297542 114656 297548 114708
rect 297600 114696 297606 114708
rect 307662 114696 307668 114708
rect 297600 114668 307668 114696
rect 297600 114656 297606 114668
rect 307662 114656 307668 114668
rect 307720 114656 307726 114708
rect 294690 114588 294696 114640
rect 294748 114628 294754 114640
rect 307570 114628 307576 114640
rect 294748 114600 307576 114628
rect 294748 114588 294754 114600
rect 307570 114588 307576 114600
rect 307628 114588 307634 114640
rect 211890 114520 211896 114572
rect 211948 114560 211954 114572
rect 213914 114560 213920 114572
rect 211948 114532 213920 114560
rect 211948 114520 211954 114532
rect 213914 114520 213920 114532
rect 213972 114520 213978 114572
rect 269758 114520 269764 114572
rect 269816 114560 269822 114572
rect 307110 114560 307116 114572
rect 269816 114532 307116 114560
rect 269816 114520 269822 114532
rect 307110 114520 307116 114532
rect 307168 114520 307174 114572
rect 252462 114452 252468 114504
rect 252520 114492 252526 114504
rect 275462 114492 275468 114504
rect 252520 114464 275468 114492
rect 252520 114452 252526 114464
rect 275462 114452 275468 114464
rect 275520 114452 275526 114504
rect 324406 114452 324412 114504
rect 324464 114492 324470 114504
rect 335446 114492 335452 114504
rect 324464 114464 335452 114492
rect 324464 114452 324470 114464
rect 335446 114452 335452 114464
rect 335504 114452 335510 114504
rect 252278 114384 252284 114436
rect 252336 114424 252342 114436
rect 256142 114424 256148 114436
rect 252336 114396 256148 114424
rect 252336 114384 252342 114396
rect 256142 114384 256148 114396
rect 256200 114384 256206 114436
rect 324314 114384 324320 114436
rect 324372 114424 324378 114436
rect 333974 114424 333980 114436
rect 324372 114396 333980 114424
rect 324372 114384 324378 114396
rect 333974 114384 333980 114396
rect 334032 114384 334038 114436
rect 251726 114316 251732 114368
rect 251784 114356 251790 114368
rect 254762 114356 254768 114368
rect 251784 114328 254768 114356
rect 251784 114316 251790 114328
rect 254762 114316 254768 114328
rect 254820 114316 254826 114368
rect 284938 113296 284944 113348
rect 284996 113336 285002 113348
rect 307570 113336 307576 113348
rect 284996 113308 307576 113336
rect 284996 113296 285002 113308
rect 307570 113296 307576 113308
rect 307628 113296 307634 113348
rect 276658 113228 276664 113280
rect 276716 113268 276722 113280
rect 307662 113268 307668 113280
rect 276716 113240 307668 113268
rect 276716 113228 276722 113240
rect 307662 113228 307668 113240
rect 307720 113228 307726 113280
rect 180242 113160 180248 113212
rect 180300 113200 180306 113212
rect 213914 113200 213920 113212
rect 180300 113172 213920 113200
rect 180300 113160 180306 113172
rect 213914 113160 213920 113172
rect 213972 113160 213978 113212
rect 260098 113160 260104 113212
rect 260156 113200 260162 113212
rect 307478 113200 307484 113212
rect 260156 113172 307484 113200
rect 260156 113160 260162 113172
rect 307478 113160 307484 113172
rect 307536 113160 307542 113212
rect 252462 113092 252468 113144
rect 252520 113132 252526 113144
rect 300394 113132 300400 113144
rect 252520 113104 300400 113132
rect 252520 113092 252526 113104
rect 300394 113092 300400 113104
rect 300452 113092 300458 113144
rect 324314 113092 324320 113144
rect 324372 113132 324378 113144
rect 339494 113132 339500 113144
rect 324372 113104 339500 113132
rect 324372 113092 324378 113104
rect 339494 113092 339500 113104
rect 339552 113092 339558 113144
rect 252094 112412 252100 112464
rect 252152 112452 252158 112464
rect 303062 112452 303068 112464
rect 252152 112424 303068 112452
rect 252152 112412 252158 112424
rect 303062 112412 303068 112424
rect 303120 112412 303126 112464
rect 252462 112276 252468 112328
rect 252520 112316 252526 112328
rect 258994 112316 259000 112328
rect 252520 112288 259000 112316
rect 252520 112276 252526 112288
rect 258994 112276 259000 112288
rect 259052 112276 259058 112328
rect 301498 111936 301504 111988
rect 301556 111976 301562 111988
rect 307662 111976 307668 111988
rect 301556 111948 307668 111976
rect 301556 111936 301562 111948
rect 307662 111936 307668 111948
rect 307720 111936 307726 111988
rect 189810 111868 189816 111920
rect 189868 111908 189874 111920
rect 214006 111908 214012 111920
rect 189868 111880 214012 111908
rect 189868 111868 189874 111880
rect 214006 111868 214012 111880
rect 214064 111868 214070 111920
rect 302970 111868 302976 111920
rect 303028 111908 303034 111920
rect 307570 111908 307576 111920
rect 303028 111880 307576 111908
rect 303028 111868 303034 111880
rect 307570 111868 307576 111880
rect 307628 111868 307634 111920
rect 170490 111800 170496 111852
rect 170548 111840 170554 111852
rect 213914 111840 213920 111852
rect 170548 111812 213920 111840
rect 170548 111800 170554 111812
rect 213914 111800 213920 111812
rect 213972 111800 213978 111852
rect 297450 111800 297456 111852
rect 297508 111840 297514 111852
rect 307662 111840 307668 111852
rect 297508 111812 307668 111840
rect 297508 111800 297514 111812
rect 307662 111800 307668 111812
rect 307720 111800 307726 111852
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 11698 111772 11704 111784
rect 3200 111744 11704 111772
rect 3200 111732 3206 111744
rect 11698 111732 11704 111744
rect 11756 111732 11762 111784
rect 168282 111732 168288 111784
rect 168340 111772 168346 111784
rect 199562 111772 199568 111784
rect 168340 111744 199568 111772
rect 168340 111732 168346 111744
rect 199562 111732 199568 111744
rect 199620 111732 199626 111784
rect 252462 111732 252468 111784
rect 252520 111772 252526 111784
rect 296162 111772 296168 111784
rect 252520 111744 296168 111772
rect 252520 111732 252526 111744
rect 296162 111732 296168 111744
rect 296220 111732 296226 111784
rect 324314 111732 324320 111784
rect 324372 111772 324378 111784
rect 340874 111772 340880 111784
rect 324372 111744 340880 111772
rect 324372 111732 324378 111744
rect 340874 111732 340880 111744
rect 340932 111732 340938 111784
rect 252370 111664 252376 111716
rect 252428 111704 252434 111716
rect 272794 111704 272800 111716
rect 252428 111676 272800 111704
rect 252428 111664 252434 111676
rect 272794 111664 272800 111676
rect 272852 111664 272858 111716
rect 304442 110576 304448 110628
rect 304500 110616 304506 110628
rect 307478 110616 307484 110628
rect 304500 110588 307484 110616
rect 304500 110576 304506 110588
rect 307478 110576 307484 110588
rect 307536 110576 307542 110628
rect 177482 110508 177488 110560
rect 177540 110548 177546 110560
rect 213914 110548 213920 110560
rect 177540 110520 213920 110548
rect 177540 110508 177546 110520
rect 213914 110508 213920 110520
rect 213972 110508 213978 110560
rect 252186 110508 252192 110560
rect 252244 110548 252250 110560
rect 256234 110548 256240 110560
rect 252244 110520 256240 110548
rect 252244 110508 252250 110520
rect 256234 110508 256240 110520
rect 256292 110508 256298 110560
rect 296254 110508 296260 110560
rect 296312 110548 296318 110560
rect 307662 110548 307668 110560
rect 296312 110520 307668 110548
rect 296312 110508 296318 110520
rect 307662 110508 307668 110520
rect 307720 110508 307726 110560
rect 166442 110440 166448 110492
rect 166500 110480 166506 110492
rect 214006 110480 214012 110492
rect 166500 110452 214012 110480
rect 166500 110440 166506 110452
rect 214006 110440 214012 110452
rect 214064 110440 214070 110492
rect 272702 110440 272708 110492
rect 272760 110480 272766 110492
rect 307570 110480 307576 110492
rect 272760 110452 307576 110480
rect 272760 110440 272766 110452
rect 307570 110440 307576 110452
rect 307628 110440 307634 110492
rect 167822 110372 167828 110424
rect 167880 110412 167886 110424
rect 177574 110412 177580 110424
rect 167880 110384 177580 110412
rect 167880 110372 167886 110384
rect 177574 110372 177580 110384
rect 177632 110372 177638 110424
rect 252370 110372 252376 110424
rect 252428 110412 252434 110424
rect 300302 110412 300308 110424
rect 252428 110384 300308 110412
rect 252428 110372 252434 110384
rect 300302 110372 300308 110384
rect 300360 110372 300366 110424
rect 324406 110372 324412 110424
rect 324464 110412 324470 110424
rect 336826 110412 336832 110424
rect 324464 110384 336832 110412
rect 324464 110372 324470 110384
rect 336826 110372 336832 110384
rect 336884 110372 336890 110424
rect 252462 110304 252468 110356
rect 252520 110344 252526 110356
rect 273990 110344 273996 110356
rect 252520 110316 273996 110344
rect 252520 110304 252526 110316
rect 273990 110304 273996 110316
rect 274048 110304 274054 110356
rect 324314 110304 324320 110356
rect 324372 110344 324378 110356
rect 332594 110344 332600 110356
rect 324372 110316 332600 110344
rect 324372 110304 324378 110316
rect 332594 110304 332600 110316
rect 332652 110304 332658 110356
rect 252278 110236 252284 110288
rect 252336 110276 252342 110288
rect 256050 110276 256056 110288
rect 252336 110248 256056 110276
rect 252336 110236 252342 110248
rect 256050 110236 256056 110248
rect 256108 110236 256114 110288
rect 301590 109148 301596 109200
rect 301648 109188 301654 109200
rect 307478 109188 307484 109200
rect 301648 109160 307484 109188
rect 301648 109148 301654 109160
rect 307478 109148 307484 109160
rect 307536 109148 307542 109200
rect 195514 109080 195520 109132
rect 195572 109120 195578 109132
rect 214006 109120 214012 109132
rect 195572 109092 214012 109120
rect 195572 109080 195578 109092
rect 214006 109080 214012 109092
rect 214064 109080 214070 109132
rect 298922 109080 298928 109132
rect 298980 109120 298986 109132
rect 307570 109120 307576 109132
rect 298980 109092 307576 109120
rect 298980 109080 298986 109092
rect 307570 109080 307576 109092
rect 307628 109080 307634 109132
rect 169018 109012 169024 109064
rect 169076 109052 169082 109064
rect 213914 109052 213920 109064
rect 169076 109024 213920 109052
rect 169076 109012 169082 109024
rect 213914 109012 213920 109024
rect 213972 109012 213978 109064
rect 275370 109012 275376 109064
rect 275428 109052 275434 109064
rect 307662 109052 307668 109064
rect 275428 109024 307668 109052
rect 275428 109012 275434 109024
rect 307662 109012 307668 109024
rect 307720 109012 307726 109064
rect 168098 108944 168104 108996
rect 168156 108984 168162 108996
rect 180334 108984 180340 108996
rect 168156 108956 180340 108984
rect 168156 108944 168162 108956
rect 180334 108944 180340 108956
rect 180392 108944 180398 108996
rect 252370 108944 252376 108996
rect 252428 108984 252434 108996
rect 301774 108984 301780 108996
rect 252428 108956 301780 108984
rect 252428 108944 252434 108956
rect 301774 108944 301780 108956
rect 301832 108944 301838 108996
rect 324314 108944 324320 108996
rect 324372 108984 324378 108996
rect 342530 108984 342536 108996
rect 324372 108956 342536 108984
rect 324372 108944 324378 108956
rect 342530 108944 342536 108956
rect 342588 108944 342594 108996
rect 252462 108876 252468 108928
rect 252520 108916 252526 108928
rect 297726 108916 297732 108928
rect 252520 108888 297732 108916
rect 252520 108876 252526 108888
rect 297726 108876 297732 108888
rect 297784 108876 297790 108928
rect 251726 108808 251732 108860
rect 251784 108848 251790 108860
rect 254670 108848 254676 108860
rect 251784 108820 254676 108848
rect 251784 108808 251790 108820
rect 254670 108808 254676 108820
rect 254728 108808 254734 108860
rect 178954 108264 178960 108316
rect 179012 108304 179018 108316
rect 214742 108304 214748 108316
rect 179012 108276 214748 108304
rect 179012 108264 179018 108276
rect 214742 108264 214748 108276
rect 214800 108264 214806 108316
rect 297634 107856 297640 107908
rect 297692 107896 297698 107908
rect 307662 107896 307668 107908
rect 297692 107868 307668 107896
rect 297692 107856 297698 107868
rect 307662 107856 307668 107868
rect 307720 107856 307726 107908
rect 300394 107720 300400 107772
rect 300452 107760 300458 107772
rect 307478 107760 307484 107772
rect 300452 107732 307484 107760
rect 300452 107720 300458 107732
rect 307478 107720 307484 107732
rect 307536 107720 307542 107772
rect 182910 107652 182916 107704
rect 182968 107692 182974 107704
rect 213914 107692 213920 107704
rect 182968 107664 213920 107692
rect 182968 107652 182974 107664
rect 213914 107652 213920 107664
rect 213972 107652 213978 107704
rect 303062 107652 303068 107704
rect 303120 107692 303126 107704
rect 307570 107692 307576 107704
rect 303120 107664 307576 107692
rect 303120 107652 303126 107664
rect 307570 107652 307576 107664
rect 307628 107652 307634 107704
rect 252370 107584 252376 107636
rect 252428 107624 252434 107636
rect 305638 107624 305644 107636
rect 252428 107596 305644 107624
rect 252428 107584 252434 107596
rect 305638 107584 305644 107596
rect 305696 107584 305702 107636
rect 252462 107516 252468 107568
rect 252520 107556 252526 107568
rect 304350 107556 304356 107568
rect 252520 107528 304356 107556
rect 252520 107516 252526 107528
rect 304350 107516 304356 107528
rect 304408 107516 304414 107568
rect 252278 107448 252284 107500
rect 252336 107488 252342 107500
rect 257338 107488 257344 107500
rect 252336 107460 257344 107488
rect 252336 107448 252342 107460
rect 257338 107448 257344 107460
rect 257396 107448 257402 107500
rect 177574 106360 177580 106412
rect 177632 106400 177638 106412
rect 213914 106400 213920 106412
rect 177632 106372 213920 106400
rect 177632 106360 177638 106372
rect 213914 106360 213920 106372
rect 213972 106360 213978 106412
rect 301774 106360 301780 106412
rect 301832 106400 301838 106412
rect 307662 106400 307668 106412
rect 301832 106372 307668 106400
rect 301832 106360 301838 106372
rect 307662 106360 307668 106372
rect 307720 106360 307726 106412
rect 167822 106292 167828 106344
rect 167880 106332 167886 106344
rect 214006 106332 214012 106344
rect 167880 106304 214012 106332
rect 167880 106292 167886 106304
rect 214006 106292 214012 106304
rect 214064 106292 214070 106344
rect 304626 106292 304632 106344
rect 304684 106332 304690 106344
rect 306742 106332 306748 106344
rect 304684 106304 306748 106332
rect 304684 106292 304690 106304
rect 306742 106292 306748 106304
rect 306800 106292 306806 106344
rect 252462 106224 252468 106276
rect 252520 106264 252526 106276
rect 261478 106264 261484 106276
rect 252520 106236 261484 106264
rect 252520 106224 252526 106236
rect 261478 106224 261484 106236
rect 261536 106224 261542 106276
rect 324314 106224 324320 106276
rect 324372 106264 324378 106276
rect 352098 106264 352104 106276
rect 324372 106236 352104 106264
rect 324372 106224 324378 106236
rect 352098 106224 352104 106236
rect 352156 106224 352162 106276
rect 251174 106156 251180 106208
rect 251232 106196 251238 106208
rect 253382 106196 253388 106208
rect 251232 106168 253388 106196
rect 251232 106156 251238 106168
rect 253382 106156 253388 106168
rect 253440 106156 253446 106208
rect 304534 105584 304540 105596
rect 258046 105556 304540 105584
rect 252370 105476 252376 105528
rect 252428 105516 252434 105528
rect 258046 105516 258074 105556
rect 304534 105544 304540 105556
rect 304592 105544 304598 105596
rect 252428 105488 258074 105516
rect 252428 105476 252434 105488
rect 258718 105000 258724 105052
rect 258776 105040 258782 105052
rect 307662 105040 307668 105052
rect 258776 105012 307668 105040
rect 258776 105000 258782 105012
rect 307662 105000 307668 105012
rect 307720 105000 307726 105052
rect 188522 104864 188528 104916
rect 188580 104904 188586 104916
rect 213914 104904 213920 104916
rect 188580 104876 213920 104904
rect 188580 104864 188586 104876
rect 213914 104864 213920 104876
rect 213972 104864 213978 104916
rect 303154 104864 303160 104916
rect 303212 104904 303218 104916
rect 307570 104904 307576 104916
rect 303212 104876 307576 104904
rect 303212 104864 303218 104876
rect 307570 104864 307576 104876
rect 307628 104864 307634 104916
rect 252462 104796 252468 104848
rect 252520 104836 252526 104848
rect 290734 104836 290740 104848
rect 252520 104808 290740 104836
rect 252520 104796 252526 104808
rect 290734 104796 290740 104808
rect 290792 104796 290798 104848
rect 173158 104116 173164 104168
rect 173216 104156 173222 104168
rect 216214 104156 216220 104168
rect 173216 104128 216220 104156
rect 173216 104116 173222 104128
rect 216214 104116 216220 104128
rect 216272 104116 216278 104168
rect 279602 104156 279608 104168
rect 252480 104128 279608 104156
rect 252480 104032 252508 104128
rect 279602 104116 279608 104128
rect 279660 104116 279666 104168
rect 252462 103980 252468 104032
rect 252520 103980 252526 104032
rect 304350 103640 304356 103692
rect 304408 103680 304414 103692
rect 307478 103680 307484 103692
rect 304408 103652 307484 103680
rect 304408 103640 304414 103652
rect 307478 103640 307484 103652
rect 307536 103640 307542 103692
rect 206554 103572 206560 103624
rect 206612 103612 206618 103624
rect 214006 103612 214012 103624
rect 206612 103584 214012 103612
rect 206612 103572 206618 103584
rect 214006 103572 214012 103584
rect 214064 103572 214070 103624
rect 290458 103572 290464 103624
rect 290516 103612 290522 103624
rect 307570 103612 307576 103624
rect 290516 103584 307576 103612
rect 290516 103572 290522 103584
rect 307570 103572 307576 103584
rect 307628 103572 307634 103624
rect 192570 103504 192576 103556
rect 192628 103544 192634 103556
rect 213914 103544 213920 103556
rect 192628 103516 213920 103544
rect 192628 103504 192634 103516
rect 213914 103504 213920 103516
rect 213972 103504 213978 103556
rect 279510 103504 279516 103556
rect 279568 103544 279574 103556
rect 307662 103544 307668 103556
rect 279568 103516 307668 103544
rect 279568 103504 279574 103516
rect 307662 103504 307668 103516
rect 307720 103504 307726 103556
rect 324498 103436 324504 103488
rect 324556 103476 324562 103488
rect 357434 103476 357440 103488
rect 324556 103448 357440 103476
rect 324556 103436 324562 103448
rect 357434 103436 357440 103448
rect 357492 103436 357498 103488
rect 324314 103300 324320 103352
rect 324372 103340 324378 103352
rect 324682 103340 324688 103352
rect 324372 103312 324688 103340
rect 324372 103300 324378 103312
rect 324682 103300 324688 103312
rect 324740 103300 324746 103352
rect 252278 103164 252284 103216
rect 252336 103204 252342 103216
rect 253290 103204 253296 103216
rect 252336 103176 253296 103204
rect 252336 103164 252342 103176
rect 253290 103164 253296 103176
rect 253348 103164 253354 103216
rect 324314 103164 324320 103216
rect 324372 103204 324378 103216
rect 327074 103204 327080 103216
rect 324372 103176 327080 103204
rect 324372 103164 324378 103176
rect 327074 103164 327080 103176
rect 327132 103164 327138 103216
rect 252186 103096 252192 103148
rect 252244 103136 252250 103148
rect 257430 103136 257436 103148
rect 252244 103108 257436 103136
rect 252244 103096 252250 103108
rect 257430 103096 257436 103108
rect 257488 103096 257494 103148
rect 289170 102280 289176 102332
rect 289228 102320 289234 102332
rect 307570 102320 307576 102332
rect 289228 102292 307576 102320
rect 289228 102280 289234 102292
rect 307570 102280 307576 102292
rect 307628 102280 307634 102332
rect 203702 102212 203708 102264
rect 203760 102252 203766 102264
rect 213914 102252 213920 102264
rect 203760 102224 213920 102252
rect 203760 102212 203766 102224
rect 213914 102212 213920 102224
rect 213972 102212 213978 102264
rect 257338 102212 257344 102264
rect 257396 102252 257402 102264
rect 307662 102252 307668 102264
rect 257396 102224 307668 102252
rect 257396 102212 257402 102224
rect 307662 102212 307668 102224
rect 307720 102212 307726 102264
rect 199562 102144 199568 102196
rect 199620 102184 199626 102196
rect 214006 102184 214012 102196
rect 199620 102156 214012 102184
rect 199620 102144 199626 102156
rect 214006 102144 214012 102156
rect 214064 102144 214070 102196
rect 253382 102144 253388 102196
rect 253440 102184 253446 102196
rect 307478 102184 307484 102196
rect 253440 102156 307484 102184
rect 253440 102144 253446 102156
rect 307478 102144 307484 102156
rect 307536 102144 307542 102196
rect 252462 102076 252468 102128
rect 252520 102116 252526 102128
rect 276750 102116 276756 102128
rect 252520 102088 276756 102116
rect 252520 102076 252526 102088
rect 276750 102076 276756 102088
rect 276808 102076 276814 102128
rect 169294 101396 169300 101448
rect 169352 101436 169358 101448
rect 214466 101436 214472 101448
rect 169352 101408 214472 101436
rect 169352 101396 169358 101408
rect 214466 101396 214472 101408
rect 214524 101396 214530 101448
rect 252186 101396 252192 101448
rect 252244 101436 252250 101448
rect 267182 101436 267188 101448
rect 252244 101408 267188 101436
rect 252244 101396 252250 101408
rect 267182 101396 267188 101408
rect 267240 101396 267246 101448
rect 267090 100920 267096 100972
rect 267148 100960 267154 100972
rect 307570 100960 307576 100972
rect 267148 100932 307576 100960
rect 267148 100920 267154 100932
rect 307570 100920 307576 100932
rect 307628 100920 307634 100972
rect 293402 100852 293408 100904
rect 293460 100892 293466 100904
rect 307662 100892 307668 100904
rect 293460 100864 307668 100892
rect 293460 100852 293466 100864
rect 307662 100852 307668 100864
rect 307720 100852 307726 100904
rect 206462 100784 206468 100836
rect 206520 100824 206526 100836
rect 214006 100824 214012 100836
rect 206520 100796 214012 100824
rect 206520 100784 206526 100796
rect 214006 100784 214012 100796
rect 214064 100784 214070 100836
rect 273990 100784 273996 100836
rect 274048 100824 274054 100836
rect 307478 100824 307484 100836
rect 274048 100796 307484 100824
rect 274048 100784 274054 100796
rect 307478 100784 307484 100796
rect 307536 100784 307542 100836
rect 173158 100716 173164 100768
rect 173216 100756 173222 100768
rect 213914 100756 213920 100768
rect 173216 100728 213920 100756
rect 173216 100716 173222 100728
rect 213914 100716 213920 100728
rect 213972 100716 213978 100768
rect 252278 100648 252284 100700
rect 252336 100688 252342 100700
rect 296346 100688 296352 100700
rect 252336 100660 296352 100688
rect 252336 100648 252342 100660
rect 296346 100648 296352 100660
rect 296404 100648 296410 100700
rect 324314 100648 324320 100700
rect 324372 100688 324378 100700
rect 331490 100688 331496 100700
rect 324372 100660 331496 100688
rect 324372 100648 324378 100660
rect 331490 100648 331496 100660
rect 331548 100648 331554 100700
rect 468478 100648 468484 100700
rect 468536 100688 468542 100700
rect 580166 100688 580172 100700
rect 468536 100660 580172 100688
rect 468536 100648 468542 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 252462 100580 252468 100632
rect 252520 100620 252526 100632
rect 294874 100620 294880 100632
rect 252520 100592 294880 100620
rect 252520 100580 252526 100592
rect 294874 100580 294880 100592
rect 294932 100580 294938 100632
rect 252370 100512 252376 100564
rect 252428 100552 252434 100564
rect 269942 100552 269948 100564
rect 252428 100524 269948 100552
rect 252428 100512 252434 100524
rect 269942 100512 269948 100524
rect 270000 100512 270006 100564
rect 300302 99492 300308 99544
rect 300360 99532 300366 99544
rect 306742 99532 306748 99544
rect 300360 99504 306748 99532
rect 300360 99492 300366 99504
rect 306742 99492 306748 99504
rect 306800 99492 306806 99544
rect 296162 99424 296168 99476
rect 296220 99464 296226 99476
rect 307662 99464 307668 99476
rect 296220 99436 307668 99464
rect 296220 99424 296226 99436
rect 307662 99424 307668 99436
rect 307720 99424 307726 99476
rect 294782 99356 294788 99408
rect 294840 99396 294846 99408
rect 307570 99396 307576 99408
rect 294840 99368 307576 99396
rect 294840 99356 294846 99368
rect 307570 99356 307576 99368
rect 307628 99356 307634 99408
rect 252462 99220 252468 99272
rect 252520 99260 252526 99272
rect 264514 99260 264520 99272
rect 252520 99232 264520 99260
rect 252520 99220 252526 99232
rect 264514 99220 264520 99232
rect 264572 99220 264578 99272
rect 252370 99152 252376 99204
rect 252428 99192 252434 99204
rect 286686 99192 286692 99204
rect 252428 99164 286692 99192
rect 252428 99152 252434 99164
rect 286686 99152 286692 99164
rect 286744 99152 286750 99204
rect 166534 98064 166540 98116
rect 166592 98104 166598 98116
rect 214006 98104 214012 98116
rect 166592 98076 214012 98104
rect 166592 98064 166598 98076
rect 214006 98064 214012 98076
rect 214064 98064 214070 98116
rect 286594 98064 286600 98116
rect 286652 98104 286658 98116
rect 307570 98104 307576 98116
rect 286652 98076 307576 98104
rect 286652 98064 286658 98076
rect 307570 98064 307576 98076
rect 307628 98064 307634 98116
rect 164878 97996 164884 98048
rect 164936 98036 164942 98048
rect 213914 98036 213920 98048
rect 164936 98008 213920 98036
rect 164936 97996 164942 98008
rect 213914 97996 213920 98008
rect 213972 97996 213978 98048
rect 261478 97996 261484 98048
rect 261536 98036 261542 98048
rect 307662 98036 307668 98048
rect 261536 98008 307668 98036
rect 261536 97996 261542 98008
rect 307662 97996 307668 98008
rect 307720 97996 307726 98048
rect 3510 97928 3516 97980
rect 3568 97968 3574 97980
rect 17218 97968 17224 97980
rect 3568 97940 17224 97968
rect 3568 97928 3574 97940
rect 17218 97928 17224 97940
rect 17276 97928 17282 97980
rect 167914 97248 167920 97300
rect 167972 97288 167978 97300
rect 214098 97288 214104 97300
rect 167972 97260 214104 97288
rect 167972 97248 167978 97260
rect 214098 97248 214104 97260
rect 214156 97248 214162 97300
rect 252462 97248 252468 97300
rect 252520 97288 252526 97300
rect 272610 97288 272616 97300
rect 252520 97260 272616 97288
rect 252520 97248 252526 97260
rect 272610 97248 272616 97260
rect 272668 97248 272674 97300
rect 291930 96772 291936 96824
rect 291988 96812 291994 96824
rect 307662 96812 307668 96824
rect 291988 96784 307668 96812
rect 291988 96772 291994 96784
rect 307662 96772 307668 96784
rect 307720 96772 307726 96824
rect 278222 96704 278228 96756
rect 278280 96744 278286 96756
rect 306926 96744 306932 96756
rect 278280 96716 306932 96744
rect 278280 96704 278286 96716
rect 306926 96704 306932 96716
rect 306984 96704 306990 96756
rect 253198 96636 253204 96688
rect 253256 96676 253262 96688
rect 307662 96676 307668 96688
rect 253256 96648 307668 96676
rect 253256 96636 253262 96648
rect 307662 96636 307668 96648
rect 307720 96636 307726 96688
rect 199470 96568 199476 96620
rect 199528 96608 199534 96620
rect 321278 96608 321284 96620
rect 199528 96580 321284 96608
rect 199528 96568 199534 96580
rect 321278 96568 321284 96580
rect 321336 96568 321342 96620
rect 286318 96500 286324 96552
rect 286376 96540 286382 96552
rect 321462 96540 321468 96552
rect 286376 96512 321468 96540
rect 286376 96500 286382 96512
rect 321462 96500 321468 96512
rect 321520 96500 321526 96552
rect 249058 95208 249064 95260
rect 249116 95248 249122 95260
rect 306926 95248 306932 95260
rect 249116 95220 306932 95248
rect 249116 95208 249122 95220
rect 306926 95208 306932 95220
rect 306984 95208 306990 95260
rect 210418 95140 210424 95192
rect 210476 95180 210482 95192
rect 324406 95180 324412 95192
rect 210476 95152 324412 95180
rect 210476 95140 210482 95152
rect 324406 95140 324412 95152
rect 324464 95140 324470 95192
rect 216122 95072 216128 95124
rect 216180 95112 216186 95124
rect 324682 95112 324688 95124
rect 216180 95084 324688 95112
rect 216180 95072 216186 95084
rect 324682 95072 324688 95084
rect 324740 95072 324746 95124
rect 59262 95004 59268 95056
rect 59320 95044 59326 95056
rect 206554 95044 206560 95056
rect 59320 95016 206560 95044
rect 59320 95004 59326 95016
rect 206554 95004 206560 95016
rect 206612 95004 206618 95056
rect 308490 95004 308496 95056
rect 308548 95044 308554 95056
rect 321554 95044 321560 95056
rect 308548 95016 321560 95044
rect 308548 95004 308554 95016
rect 321554 95004 321560 95016
rect 321612 95004 321618 95056
rect 162854 94528 162860 94580
rect 162912 94568 162918 94580
rect 203610 94568 203616 94580
rect 162912 94540 203616 94568
rect 162912 94528 162918 94540
rect 203610 94528 203616 94540
rect 203668 94528 203674 94580
rect 122834 94460 122840 94512
rect 122892 94500 122898 94512
rect 214650 94500 214656 94512
rect 122892 94472 214656 94500
rect 122892 94460 122898 94472
rect 214650 94460 214656 94472
rect 214708 94460 214714 94512
rect 151722 93916 151728 93968
rect 151780 93956 151786 93968
rect 178862 93956 178868 93968
rect 151780 93928 178868 93956
rect 151780 93916 151786 93928
rect 178862 93916 178868 93928
rect 178920 93916 178926 93968
rect 129366 93848 129372 93900
rect 129424 93888 129430 93900
rect 167730 93888 167736 93900
rect 129424 93860 167736 93888
rect 129424 93848 129430 93860
rect 167730 93848 167736 93860
rect 167788 93848 167794 93900
rect 151722 93440 151728 93492
rect 151780 93480 151786 93492
rect 175918 93480 175924 93492
rect 151780 93452 175924 93480
rect 151780 93440 151786 93452
rect 175918 93440 175924 93452
rect 175976 93440 175982 93492
rect 135714 93372 135720 93424
rect 135772 93412 135778 93424
rect 167638 93412 167644 93424
rect 135772 93384 167644 93412
rect 135772 93372 135778 93384
rect 167638 93372 167644 93384
rect 167696 93372 167702 93424
rect 120626 93304 120632 93356
rect 120684 93344 120690 93356
rect 170582 93344 170588 93356
rect 120684 93316 170588 93344
rect 120684 93304 120690 93316
rect 170582 93304 170588 93316
rect 170640 93304 170646 93356
rect 115474 93236 115480 93288
rect 115532 93276 115538 93288
rect 166258 93276 166264 93288
rect 115532 93248 166264 93276
rect 115532 93236 115538 93248
rect 166258 93236 166264 93248
rect 166316 93236 166322 93288
rect 85666 93168 85672 93220
rect 85724 93208 85730 93220
rect 164878 93208 164884 93220
rect 85724 93180 164884 93208
rect 85724 93168 85730 93180
rect 164878 93168 164884 93180
rect 164936 93168 164942 93220
rect 126606 93100 126612 93152
rect 126664 93140 126670 93152
rect 214834 93140 214840 93152
rect 126664 93112 214840 93140
rect 126664 93100 126670 93112
rect 214834 93100 214840 93112
rect 214892 93100 214898 93152
rect 238018 93100 238024 93152
rect 238076 93140 238082 93152
rect 251174 93140 251180 93152
rect 238076 93112 251180 93140
rect 238076 93100 238082 93112
rect 251174 93100 251180 93112
rect 251232 93100 251238 93152
rect 74810 92420 74816 92472
rect 74868 92460 74874 92472
rect 214742 92460 214748 92472
rect 74868 92432 214748 92460
rect 74868 92420 74874 92432
rect 214742 92420 214748 92432
rect 214800 92420 214806 92472
rect 88978 92352 88984 92404
rect 89036 92392 89042 92404
rect 167914 92392 167920 92404
rect 89036 92364 167920 92392
rect 89036 92352 89042 92364
rect 167914 92352 167920 92364
rect 167972 92352 167978 92404
rect 95050 92284 95056 92336
rect 95108 92324 95114 92336
rect 122834 92324 122840 92336
rect 95108 92296 122840 92324
rect 95108 92284 95114 92296
rect 122834 92284 122840 92296
rect 122892 92284 122898 92336
rect 134426 92284 134432 92336
rect 134484 92324 134490 92336
rect 210602 92324 210608 92336
rect 134484 92296 210608 92324
rect 134484 92284 134490 92296
rect 210602 92284 210608 92296
rect 210660 92284 210666 92336
rect 105538 92216 105544 92268
rect 105596 92256 105602 92268
rect 126606 92256 126612 92268
rect 105596 92228 126612 92256
rect 105596 92216 105602 92228
rect 126606 92216 126612 92228
rect 126664 92216 126670 92268
rect 126698 92216 126704 92268
rect 126756 92256 126762 92268
rect 202230 92256 202236 92268
rect 126756 92228 202236 92256
rect 126756 92216 126762 92228
rect 202230 92216 202236 92228
rect 202288 92216 202294 92268
rect 116762 92148 116768 92200
rect 116820 92188 116826 92200
rect 169294 92188 169300 92200
rect 116820 92160 169300 92188
rect 116820 92148 116826 92160
rect 169294 92148 169300 92160
rect 169352 92148 169358 92200
rect 128170 92080 128176 92132
rect 128228 92120 128234 92132
rect 173434 92120 173440 92132
rect 128228 92092 173440 92120
rect 128228 92080 128234 92092
rect 173434 92080 173440 92092
rect 173492 92080 173498 92132
rect 178678 91740 178684 91792
rect 178736 91780 178742 91792
rect 307294 91780 307300 91792
rect 178736 91752 307300 91780
rect 178736 91740 178742 91752
rect 307294 91740 307300 91752
rect 307352 91740 307358 91792
rect 102042 91060 102048 91112
rect 102100 91100 102106 91112
rect 118694 91100 118700 91112
rect 102100 91072 118700 91100
rect 102100 91060 102106 91072
rect 118694 91060 118700 91072
rect 118752 91060 118758 91112
rect 67358 90992 67364 91044
rect 67416 91032 67422 91044
rect 203702 91032 203708 91044
rect 67416 91004 203708 91032
rect 67416 90992 67422 91004
rect 203702 90992 203708 91004
rect 203760 90992 203766 91044
rect 62022 90924 62028 90976
rect 62080 90964 62086 90976
rect 192570 90964 192576 90976
rect 62080 90936 192576 90964
rect 62080 90924 62086 90936
rect 192570 90924 192576 90936
rect 192628 90924 192634 90976
rect 106642 90856 106648 90908
rect 106700 90896 106706 90908
rect 173342 90896 173348 90908
rect 106700 90868 173348 90896
rect 106700 90856 106706 90868
rect 173342 90856 173348 90868
rect 173400 90856 173406 90908
rect 110322 90788 110328 90840
rect 110380 90828 110386 90840
rect 170674 90828 170680 90840
rect 110380 90800 170680 90828
rect 110380 90788 110386 90800
rect 170674 90788 170680 90800
rect 170732 90788 170738 90840
rect 124030 90720 124036 90772
rect 124088 90760 124094 90772
rect 169202 90760 169208 90772
rect 124088 90732 169208 90760
rect 124088 90720 124094 90732
rect 169202 90720 169208 90732
rect 169260 90720 169266 90772
rect 151722 90652 151728 90704
rect 151780 90692 151786 90704
rect 177298 90692 177304 90704
rect 151780 90664 177304 90692
rect 151780 90652 151786 90664
rect 177298 90652 177304 90664
rect 177356 90652 177362 90704
rect 115566 89632 115572 89684
rect 115624 89672 115630 89684
rect 213362 89672 213368 89684
rect 115624 89644 213368 89672
rect 115624 89632 115630 89644
rect 213362 89632 213368 89644
rect 213420 89632 213426 89684
rect 113818 89564 113824 89616
rect 113876 89604 113882 89616
rect 185670 89604 185676 89616
rect 113876 89576 185676 89604
rect 113876 89564 113882 89576
rect 185670 89564 185676 89576
rect 185728 89564 185734 89616
rect 118694 89496 118700 89548
rect 118752 89536 118758 89548
rect 189810 89536 189816 89548
rect 118752 89508 189816 89536
rect 118752 89496 118758 89508
rect 189810 89496 189816 89508
rect 189868 89496 189874 89548
rect 126882 89428 126888 89480
rect 126940 89468 126946 89480
rect 176102 89468 176108 89480
rect 126940 89440 176108 89468
rect 126940 89428 126946 89440
rect 176102 89428 176108 89440
rect 176160 89428 176166 89480
rect 125410 89360 125416 89412
rect 125468 89400 125474 89412
rect 171778 89400 171784 89412
rect 125468 89372 171784 89400
rect 125468 89360 125474 89372
rect 171778 89360 171784 89372
rect 171836 89360 171842 89412
rect 153010 89292 153016 89344
rect 153068 89332 153074 89344
rect 184290 89332 184296 89344
rect 153068 89304 184296 89332
rect 153068 89292 153074 89304
rect 184290 89292 184296 89304
rect 184348 89292 184354 89344
rect 188338 88952 188344 89004
rect 188396 88992 188402 89004
rect 324314 88992 324320 89004
rect 188396 88964 324320 88992
rect 188396 88952 188402 88964
rect 324314 88952 324320 88964
rect 324372 88952 324378 89004
rect 107194 88272 107200 88324
rect 107252 88312 107258 88324
rect 211890 88312 211896 88324
rect 107252 88284 211896 88312
rect 107252 88272 107258 88284
rect 211890 88272 211896 88284
rect 211948 88272 211954 88324
rect 90726 88204 90732 88256
rect 90784 88244 90790 88256
rect 188522 88244 188528 88256
rect 90784 88216 188528 88244
rect 90784 88204 90790 88216
rect 188522 88204 188528 88216
rect 188580 88204 188586 88256
rect 100202 88136 100208 88188
rect 100260 88176 100266 88188
rect 166442 88176 166448 88188
rect 100260 88148 166448 88176
rect 100260 88136 100266 88148
rect 166442 88136 166448 88148
rect 166500 88136 166506 88188
rect 118234 88068 118240 88120
rect 118292 88108 118298 88120
rect 177390 88108 177396 88120
rect 118292 88080 177396 88108
rect 118292 88068 118298 88080
rect 177390 88068 177396 88080
rect 177448 88068 177454 88120
rect 132402 88000 132408 88052
rect 132460 88040 132466 88052
rect 174630 88040 174636 88052
rect 132460 88012 174636 88040
rect 132460 88000 132466 88012
rect 174630 88000 174636 88012
rect 174688 88000 174694 88052
rect 188338 87592 188344 87644
rect 188396 87632 188402 87644
rect 307202 87632 307208 87644
rect 188396 87604 307208 87632
rect 188396 87592 188402 87604
rect 307202 87592 307208 87604
rect 307260 87592 307266 87644
rect 67634 86912 67640 86964
rect 67692 86952 67698 86964
rect 214558 86952 214564 86964
rect 67692 86924 214564 86952
rect 67692 86912 67698 86924
rect 214558 86912 214564 86924
rect 214616 86912 214622 86964
rect 97074 86844 97080 86896
rect 97132 86884 97138 86896
rect 198090 86884 198096 86896
rect 97132 86856 198096 86884
rect 97132 86844 97138 86856
rect 198090 86844 198096 86856
rect 198148 86844 198154 86896
rect 108482 86776 108488 86828
rect 108540 86816 108546 86828
rect 181530 86816 181536 86828
rect 108540 86788 181536 86816
rect 108540 86776 108546 86788
rect 181530 86776 181536 86788
rect 181588 86776 181594 86828
rect 117130 86708 117136 86760
rect 117188 86748 117194 86760
rect 166350 86748 166356 86760
rect 117188 86720 166356 86748
rect 117188 86708 117194 86720
rect 166350 86708 166356 86720
rect 166408 86708 166414 86760
rect 126698 86640 126704 86692
rect 126756 86680 126762 86692
rect 173250 86680 173256 86692
rect 126756 86652 173256 86680
rect 126756 86640 126762 86652
rect 173250 86640 173256 86652
rect 173308 86640 173314 86692
rect 202138 86232 202144 86284
rect 202196 86272 202202 86284
rect 307754 86272 307760 86284
rect 202196 86244 307760 86272
rect 202196 86232 202202 86244
rect 307754 86232 307760 86244
rect 307812 86232 307818 86284
rect 3510 85484 3516 85536
rect 3568 85524 3574 85536
rect 54478 85524 54484 85536
rect 3568 85496 54484 85524
rect 3568 85484 3574 85496
rect 54478 85484 54484 85496
rect 54536 85484 54542 85536
rect 102962 85484 102968 85536
rect 103020 85524 103026 85536
rect 213454 85524 213460 85536
rect 103020 85496 213460 85524
rect 103020 85484 103026 85496
rect 213454 85484 213460 85496
rect 213512 85484 213518 85536
rect 108206 85416 108212 85468
rect 108264 85456 108270 85468
rect 202322 85456 202328 85468
rect 108264 85428 202328 85456
rect 108264 85416 108270 85428
rect 202322 85416 202328 85428
rect 202380 85416 202386 85468
rect 109586 85348 109592 85400
rect 109644 85388 109650 85400
rect 181438 85388 181444 85400
rect 109644 85360 181444 85388
rect 109644 85348 109650 85360
rect 181438 85348 181444 85360
rect 181496 85348 181502 85400
rect 122834 85280 122840 85332
rect 122892 85320 122898 85332
rect 187142 85320 187148 85332
rect 122892 85292 187148 85320
rect 122892 85280 122898 85292
rect 187142 85280 187148 85292
rect 187200 85280 187206 85332
rect 112530 85212 112536 85264
rect 112588 85252 112594 85264
rect 170398 85252 170404 85264
rect 112588 85224 170404 85252
rect 112588 85212 112594 85224
rect 170398 85212 170404 85224
rect 170456 85212 170462 85264
rect 133230 85144 133236 85196
rect 133288 85184 133294 85196
rect 174538 85184 174544 85196
rect 133288 85156 174544 85184
rect 133288 85144 133294 85156
rect 174538 85144 174544 85156
rect 174596 85144 174602 85196
rect 206278 84804 206284 84856
rect 206336 84844 206342 84856
rect 324406 84844 324412 84856
rect 206336 84816 324412 84844
rect 206336 84804 206342 84816
rect 324406 84804 324412 84816
rect 324464 84804 324470 84856
rect 67542 84124 67548 84176
rect 67600 84164 67606 84176
rect 206462 84164 206468 84176
rect 67600 84136 206468 84164
rect 67600 84124 67606 84136
rect 206462 84124 206468 84136
rect 206520 84124 206526 84176
rect 115842 84056 115848 84108
rect 115900 84096 115906 84108
rect 188430 84096 188436 84108
rect 115900 84068 188436 84096
rect 115900 84056 115906 84068
rect 188430 84056 188436 84068
rect 188488 84056 188494 84108
rect 96522 83988 96528 84040
rect 96580 84028 96586 84040
rect 169018 84028 169024 84040
rect 96580 84000 169024 84028
rect 96580 83988 96586 84000
rect 169018 83988 169024 84000
rect 169076 83988 169082 84040
rect 111702 83920 111708 83972
rect 111760 83960 111766 83972
rect 174722 83960 174728 83972
rect 111760 83932 174728 83960
rect 111760 83920 111766 83932
rect 174722 83920 174728 83932
rect 174780 83920 174786 83972
rect 196618 83444 196624 83496
rect 196676 83484 196682 83496
rect 314654 83484 314660 83496
rect 196676 83456 314660 83484
rect 196676 83444 196682 83456
rect 314654 83444 314660 83456
rect 314712 83444 314718 83496
rect 110138 82764 110144 82816
rect 110196 82804 110202 82816
rect 198182 82804 198188 82816
rect 110196 82776 198188 82804
rect 110196 82764 110202 82776
rect 198182 82764 198188 82776
rect 198240 82764 198246 82816
rect 124122 82696 124128 82748
rect 124180 82736 124186 82748
rect 210510 82736 210516 82748
rect 124180 82708 210516 82736
rect 124180 82696 124186 82708
rect 210510 82696 210516 82708
rect 210568 82696 210574 82748
rect 99190 82628 99196 82680
rect 99248 82668 99254 82680
rect 177482 82668 177488 82680
rect 99248 82640 177488 82668
rect 99248 82628 99254 82640
rect 177482 82628 177488 82640
rect 177540 82628 177546 82680
rect 101950 82560 101956 82612
rect 102008 82600 102014 82612
rect 171962 82600 171968 82612
rect 102008 82572 171968 82600
rect 102008 82560 102014 82572
rect 171962 82560 171968 82572
rect 172020 82560 172026 82612
rect 122650 82492 122656 82544
rect 122708 82532 122714 82544
rect 169110 82532 169116 82544
rect 122708 82504 169116 82532
rect 122708 82492 122714 82504
rect 169110 82492 169116 82504
rect 169168 82492 169174 82544
rect 206370 82084 206376 82136
rect 206428 82124 206434 82136
rect 329834 82124 329840 82136
rect 206428 82096 329840 82124
rect 206428 82084 206434 82096
rect 329834 82084 329840 82096
rect 329892 82084 329898 82136
rect 92382 81336 92388 81388
rect 92440 81376 92446 81388
rect 177574 81376 177580 81388
rect 92440 81348 177580 81376
rect 92440 81336 92446 81348
rect 177574 81336 177580 81348
rect 177632 81336 177638 81388
rect 125502 81268 125508 81320
rect 125560 81308 125566 81320
rect 207750 81308 207756 81320
rect 125560 81280 207756 81308
rect 125560 81268 125566 81280
rect 207750 81268 207756 81280
rect 207808 81268 207814 81320
rect 100662 81200 100668 81252
rect 100720 81240 100726 81252
rect 170490 81240 170496 81252
rect 100720 81212 170496 81240
rect 100720 81200 100726 81212
rect 170490 81200 170496 81212
rect 170548 81200 170554 81252
rect 104710 81132 104716 81184
rect 104768 81172 104774 81184
rect 171870 81172 171876 81184
rect 104768 81144 171876 81172
rect 104768 81132 104774 81144
rect 171870 81132 171876 81144
rect 171928 81132 171934 81184
rect 131022 81064 131028 81116
rect 131080 81104 131086 81116
rect 184198 81104 184204 81116
rect 131080 81076 184204 81104
rect 131080 81064 131086 81076
rect 184198 81064 184204 81076
rect 184256 81064 184262 81116
rect 209038 80656 209044 80708
rect 209096 80696 209102 80708
rect 325694 80696 325700 80708
rect 209096 80668 325700 80696
rect 209096 80656 209102 80668
rect 325694 80656 325700 80668
rect 325752 80656 325758 80708
rect 119982 79976 119988 80028
rect 120040 80016 120046 80028
rect 209222 80016 209228 80028
rect 120040 79988 209228 80016
rect 120040 79976 120046 79988
rect 209222 79976 209228 79988
rect 209280 79976 209286 80028
rect 95142 79908 95148 79960
rect 95200 79948 95206 79960
rect 182910 79948 182916 79960
rect 95200 79920 182916 79948
rect 95200 79908 95206 79920
rect 182910 79908 182916 79920
rect 182968 79908 182974 79960
rect 86862 79840 86868 79892
rect 86920 79880 86926 79892
rect 166534 79880 166540 79892
rect 86920 79852 166540 79880
rect 86920 79840 86926 79852
rect 166534 79840 166540 79852
rect 166592 79840 166598 79892
rect 118602 79772 118608 79824
rect 118660 79812 118666 79824
rect 196710 79812 196716 79824
rect 118660 79784 196716 79812
rect 118660 79772 118666 79784
rect 196710 79772 196716 79784
rect 196768 79772 196774 79824
rect 97902 78616 97908 78668
rect 97960 78656 97966 78668
rect 195514 78656 195520 78668
rect 97960 78628 195520 78656
rect 97960 78616 97966 78628
rect 195514 78616 195520 78628
rect 195572 78616 195578 78668
rect 122742 78548 122748 78600
rect 122800 78588 122806 78600
rect 213270 78588 213276 78600
rect 122800 78560 213276 78588
rect 122800 78548 122806 78560
rect 213270 78548 213276 78560
rect 213328 78548 213334 78600
rect 93762 78480 93768 78532
rect 93820 78520 93826 78532
rect 167822 78520 167828 78532
rect 93820 78492 167828 78520
rect 93820 78480 93826 78492
rect 167822 78480 167828 78492
rect 167880 78480 167886 78532
rect 101858 78412 101864 78464
rect 101916 78452 101922 78464
rect 176010 78452 176016 78464
rect 101916 78424 176016 78452
rect 101916 78412 101922 78424
rect 176010 78412 176016 78424
rect 176068 78412 176074 78464
rect 211798 78004 211804 78056
rect 211856 78044 211862 78056
rect 260834 78044 260840 78056
rect 211856 78016 260840 78044
rect 211856 78004 211862 78016
rect 260834 78004 260840 78016
rect 260892 78004 260898 78056
rect 280798 78004 280804 78056
rect 280856 78044 280862 78056
rect 316034 78044 316040 78056
rect 280856 78016 316040 78044
rect 280856 78004 280862 78016
rect 316034 78004 316040 78016
rect 316092 78004 316098 78056
rect 180058 77936 180064 77988
rect 180116 77976 180122 77988
rect 321554 77976 321560 77988
rect 180116 77948 321560 77976
rect 180116 77936 180122 77948
rect 321554 77936 321560 77948
rect 321612 77936 321618 77988
rect 85482 77188 85488 77240
rect 85540 77228 85546 77240
rect 173158 77228 173164 77240
rect 85540 77200 173164 77228
rect 85540 77188 85546 77200
rect 173158 77188 173164 77200
rect 173216 77188 173222 77240
rect 121362 77120 121368 77172
rect 121420 77160 121426 77172
rect 207658 77160 207664 77172
rect 121420 77132 207664 77160
rect 121420 77120 121426 77132
rect 207658 77120 207664 77132
rect 207716 77120 207722 77172
rect 114462 77052 114468 77104
rect 114520 77092 114526 77104
rect 178770 77092 178776 77104
rect 114520 77064 178776 77092
rect 114520 77052 114526 77064
rect 178770 77052 178776 77064
rect 178828 77052 178834 77104
rect 92474 76508 92480 76560
rect 92532 76548 92538 76560
rect 300210 76548 300216 76560
rect 92532 76520 300216 76548
rect 92532 76508 92538 76520
rect 300210 76508 300216 76520
rect 300268 76508 300274 76560
rect 104802 75828 104808 75880
rect 104860 75868 104866 75880
rect 180242 75868 180248 75880
rect 104860 75840 180248 75868
rect 104860 75828 104866 75840
rect 180242 75828 180248 75840
rect 180300 75828 180306 75880
rect 95234 75216 95240 75268
rect 95292 75256 95298 75268
rect 265710 75256 265716 75268
rect 95292 75228 265716 75256
rect 95292 75216 95298 75228
rect 265710 75216 265716 75228
rect 265768 75216 265774 75268
rect 69014 75148 69020 75200
rect 69072 75188 69078 75200
rect 303154 75188 303160 75200
rect 69072 75160 303160 75188
rect 69072 75148 69078 75160
rect 303154 75148 303160 75160
rect 303212 75148 303218 75200
rect 122834 73924 122840 73976
rect 122892 73964 122898 73976
rect 254578 73964 254584 73976
rect 122892 73936 254584 73964
rect 122892 73924 122898 73936
rect 254578 73924 254584 73936
rect 254636 73924 254642 73976
rect 99374 73856 99380 73908
rect 99432 73896 99438 73908
rect 285030 73896 285036 73908
rect 99432 73868 285036 73896
rect 99432 73856 99438 73868
rect 285030 73856 285036 73868
rect 285088 73856 285094 73908
rect 71774 73788 71780 73840
rect 71832 73828 71838 73840
rect 305914 73828 305920 73840
rect 71832 73800 305920 73828
rect 71832 73788 71838 73800
rect 305914 73788 305920 73800
rect 305972 73788 305978 73840
rect 115934 72564 115940 72616
rect 115992 72604 115998 72616
rect 255958 72604 255964 72616
rect 115992 72576 255964 72604
rect 115992 72564 115998 72576
rect 255958 72564 255964 72576
rect 256016 72564 256022 72616
rect 84194 72496 84200 72548
rect 84252 72536 84258 72548
rect 271230 72536 271236 72548
rect 84252 72508 271236 72536
rect 84252 72496 84258 72508
rect 271230 72496 271236 72508
rect 271288 72496 271294 72548
rect 67634 72428 67640 72480
rect 67692 72468 67698 72480
rect 273898 72468 273904 72480
rect 67692 72440 273904 72468
rect 67692 72428 67698 72440
rect 273898 72428 273904 72440
rect 273956 72428 273962 72480
rect 97994 71068 98000 71120
rect 98052 71108 98058 71120
rect 301682 71108 301688 71120
rect 98052 71080 301688 71108
rect 98052 71068 98058 71080
rect 301682 71068 301688 71080
rect 301740 71068 301746 71120
rect 46934 71000 46940 71052
rect 46992 71040 46998 71052
rect 253382 71040 253388 71052
rect 46992 71012 253388 71040
rect 46992 71000 46998 71012
rect 253382 71000 253388 71012
rect 253440 71000 253446 71052
rect 110414 69708 110420 69760
rect 110472 69748 110478 69760
rect 292022 69748 292028 69760
rect 110472 69720 292028 69748
rect 110472 69708 110478 69720
rect 292022 69708 292028 69720
rect 292080 69708 292086 69760
rect 75914 69640 75920 69692
rect 75972 69680 75978 69692
rect 304626 69680 304632 69692
rect 75972 69652 304632 69680
rect 75972 69640 75978 69652
rect 304626 69640 304632 69652
rect 304684 69640 304690 69692
rect 113174 68416 113180 68468
rect 113232 68456 113238 68468
rect 294598 68456 294604 68468
rect 113232 68428 294604 68456
rect 113232 68416 113238 68428
rect 294598 68416 294604 68428
rect 294656 68416 294662 68468
rect 78674 68348 78680 68400
rect 78732 68388 78738 68400
rect 301774 68388 301780 68400
rect 78732 68360 301780 68388
rect 78732 68348 78738 68360
rect 301774 68348 301780 68360
rect 301832 68348 301838 68400
rect 4154 68280 4160 68332
rect 4212 68320 4218 68332
rect 249058 68320 249064 68332
rect 4212 68292 249064 68320
rect 4212 68280 4218 68292
rect 249058 68280 249064 68292
rect 249116 68280 249122 68332
rect 82814 66920 82820 66972
rect 82872 66960 82878 66972
rect 300394 66960 300400 66972
rect 82872 66932 300400 66960
rect 82872 66920 82878 66932
rect 300394 66920 300400 66932
rect 300452 66920 300458 66972
rect 13814 66852 13820 66904
rect 13872 66892 13878 66904
rect 289354 66892 289360 66904
rect 13872 66864 289360 66892
rect 13872 66852 13878 66864
rect 289354 66852 289360 66864
rect 289412 66852 289418 66904
rect 85574 65560 85580 65612
rect 85632 65600 85638 65612
rect 305822 65600 305828 65612
rect 85632 65572 305828 65600
rect 85632 65560 85638 65572
rect 305822 65560 305828 65572
rect 305880 65560 305886 65612
rect 60734 65492 60740 65544
rect 60792 65532 60798 65544
rect 286502 65532 286508 65544
rect 60792 65504 286508 65532
rect 60792 65492 60798 65504
rect 286502 65492 286508 65504
rect 286560 65492 286566 65544
rect 89714 64132 89720 64184
rect 89772 64172 89778 64184
rect 303062 64172 303068 64184
rect 89772 64144 303068 64172
rect 89772 64132 89778 64144
rect 303062 64132 303068 64144
rect 303120 64132 303126 64184
rect 93854 62772 93860 62824
rect 93912 62812 93918 62824
rect 297634 62812 297640 62824
rect 93912 62784 297640 62812
rect 93912 62772 93918 62784
rect 297634 62772 297640 62784
rect 297692 62772 297698 62824
rect 96614 61412 96620 61464
rect 96672 61452 96678 61464
rect 275370 61452 275376 61464
rect 96672 61424 275376 61452
rect 96672 61412 96678 61424
rect 275370 61412 275376 61424
rect 275428 61412 275434 61464
rect 278038 61412 278044 61464
rect 278096 61452 278102 61464
rect 316126 61452 316132 61464
rect 278096 61424 316132 61452
rect 278096 61412 278102 61424
rect 316126 61412 316132 61424
rect 316184 61412 316190 61464
rect 44174 61344 44180 61396
rect 44232 61384 44238 61396
rect 282362 61384 282368 61396
rect 44232 61356 282368 61384
rect 44232 61344 44238 61356
rect 282362 61344 282368 61356
rect 282420 61344 282426 61396
rect 185578 60052 185584 60104
rect 185636 60092 185642 60104
rect 313274 60092 313280 60104
rect 185636 60064 313280 60092
rect 185636 60052 185642 60064
rect 313274 60052 313280 60064
rect 313332 60052 313338 60104
rect 12434 59984 12440 60036
rect 12492 60024 12498 60036
rect 276658 60024 276664 60036
rect 12492 59996 276664 60024
rect 12492 59984 12498 59996
rect 276658 59984 276664 59996
rect 276716 59984 276722 60036
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 53098 59344 53104 59356
rect 3108 59316 53104 59344
rect 3108 59304 3114 59316
rect 53098 59304 53104 59316
rect 53156 59304 53162 59356
rect 100754 58692 100760 58744
rect 100812 58732 100818 58744
rect 298922 58732 298928 58744
rect 100812 58704 298928 58732
rect 100812 58692 100818 58704
rect 298922 58692 298928 58704
rect 298980 58692 298986 58744
rect 52454 58624 52460 58676
rect 52512 58664 52518 58676
rect 290642 58664 290648 58676
rect 52512 58636 290648 58664
rect 52512 58624 52518 58636
rect 290642 58624 290648 58636
rect 290700 58624 290706 58676
rect 103514 57264 103520 57316
rect 103572 57304 103578 57316
rect 301590 57304 301596 57316
rect 103572 57276 301596 57304
rect 103572 57264 103578 57276
rect 301590 57264 301596 57276
rect 301648 57264 301654 57316
rect 37274 57196 37280 57248
rect 37332 57236 37338 57248
rect 269758 57236 269764 57248
rect 37332 57208 269764 57236
rect 37332 57196 37338 57208
rect 269758 57196 269764 57208
rect 269816 57196 269822 57248
rect 107654 55904 107660 55956
rect 107712 55944 107718 55956
rect 296254 55944 296260 55956
rect 107712 55916 296260 55944
rect 107712 55904 107718 55916
rect 296254 55904 296260 55916
rect 296312 55904 296318 55956
rect 34514 55836 34520 55888
rect 34572 55876 34578 55888
rect 294690 55876 294696 55888
rect 34572 55848 294696 55876
rect 34572 55836 34578 55848
rect 294690 55836 294696 55848
rect 294748 55836 294754 55888
rect 110506 54544 110512 54596
rect 110564 54584 110570 54596
rect 304442 54584 304448 54596
rect 110564 54556 304448 54584
rect 110564 54544 110570 54556
rect 304442 54544 304448 54556
rect 304500 54544 304506 54596
rect 30374 54476 30380 54528
rect 30432 54516 30438 54528
rect 297542 54516 297548 54528
rect 30432 54488 297548 54516
rect 30432 54476 30438 54488
rect 297542 54476 297548 54488
rect 297600 54476 297606 54528
rect 114554 53048 114560 53100
rect 114612 53088 114618 53100
rect 272702 53088 272708 53100
rect 114612 53060 272708 53088
rect 114612 53048 114618 53060
rect 272702 53048 272708 53060
rect 272760 53048 272766 53100
rect 124214 51756 124220 51808
rect 124272 51796 124278 51808
rect 282270 51796 282276 51808
rect 124272 51768 282276 51796
rect 124272 51756 124278 51768
rect 282270 51756 282276 51768
rect 282328 51756 282334 51808
rect 16574 51688 16580 51740
rect 16632 51728 16638 51740
rect 300302 51728 300308 51740
rect 16632 51700 300308 51728
rect 16632 51688 16638 51700
rect 300302 51688 300308 51700
rect 300360 51688 300366 51740
rect 81434 50396 81440 50448
rect 81492 50436 81498 50448
rect 293218 50436 293224 50448
rect 81492 50408 293224 50436
rect 81492 50396 81498 50408
rect 293218 50396 293224 50408
rect 293276 50396 293282 50448
rect 27614 50328 27620 50380
rect 27672 50368 27678 50380
rect 260098 50368 260104 50380
rect 27672 50340 260104 50368
rect 27672 50328 27678 50340
rect 260098 50328 260104 50340
rect 260156 50328 260162 50380
rect 106274 49104 106280 49156
rect 106332 49144 106338 49156
rect 250530 49144 250536 49156
rect 106332 49116 250536 49144
rect 106332 49104 106338 49116
rect 250530 49104 250536 49116
rect 250588 49104 250594 49156
rect 121454 49036 121460 49088
rect 121512 49076 121518 49088
rect 302970 49076 302976 49088
rect 121512 49048 302976 49076
rect 121512 49036 121518 49048
rect 302970 49036 302976 49048
rect 303028 49036 303034 49088
rect 17954 48968 17960 49020
rect 18012 49008 18018 49020
rect 284938 49008 284944 49020
rect 18012 48980 284944 49008
rect 18012 48968 18018 48980
rect 284938 48968 284944 48980
rect 284996 48968 285002 49020
rect 31754 47608 31760 47660
rect 31812 47648 31818 47660
rect 290550 47648 290556 47660
rect 31812 47620 290556 47648
rect 31812 47608 31818 47620
rect 290550 47608 290556 47620
rect 290608 47608 290614 47660
rect 20714 47540 20720 47592
rect 20772 47580 20778 47592
rect 294782 47580 294788 47592
rect 20772 47552 294788 47580
rect 20772 47540 20778 47552
rect 294782 47540 294788 47552
rect 294840 47540 294846 47592
rect 180150 46860 180156 46912
rect 180208 46900 180214 46912
rect 580166 46900 580172 46912
rect 180208 46872 580172 46900
rect 180208 46860 180214 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 73154 46248 73160 46300
rect 73212 46288 73218 46300
rect 262858 46288 262864 46300
rect 73212 46260 262864 46288
rect 73212 46248 73218 46260
rect 262858 46248 262864 46260
rect 262916 46248 262922 46300
rect 93946 46180 93952 46232
rect 94004 46220 94010 46232
rect 293310 46220 293316 46232
rect 94004 46192 293316 46220
rect 94004 46180 94010 46192
rect 293310 46180 293316 46192
rect 293368 46180 293374 46232
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 15838 45540 15844 45552
rect 3476 45512 15844 45540
rect 3476 45500 3482 45512
rect 15838 45500 15844 45512
rect 15896 45500 15902 45552
rect 35894 44888 35900 44940
rect 35952 44928 35958 44940
rect 271138 44928 271144 44940
rect 35952 44900 271144 44928
rect 35952 44888 35958 44900
rect 271138 44888 271144 44900
rect 271196 44888 271202 44940
rect 26234 44820 26240 44872
rect 26292 44860 26298 44872
rect 293402 44860 293408 44872
rect 26292 44832 293408 44860
rect 26292 44820 26298 44832
rect 293402 44820 293408 44832
rect 293460 44820 293466 44872
rect 88334 43460 88340 43512
rect 88392 43500 88398 43512
rect 289262 43500 289268 43512
rect 88392 43472 289268 43500
rect 88392 43460 88398 43472
rect 289262 43460 289268 43472
rect 289320 43460 289326 43512
rect 28994 43392 29000 43444
rect 29052 43432 29058 43444
rect 273990 43432 273996 43444
rect 29052 43404 273996 43432
rect 29052 43392 29058 43404
rect 273990 43392 273996 43404
rect 274048 43392 274054 43444
rect 27706 42100 27712 42152
rect 27764 42140 27770 42152
rect 280982 42140 280988 42152
rect 27764 42112 280988 42140
rect 27764 42100 27770 42112
rect 280982 42100 280988 42112
rect 281040 42100 281046 42152
rect 33134 42032 33140 42084
rect 33192 42072 33198 42084
rect 305730 42072 305736 42084
rect 33192 42044 305736 42072
rect 33192 42032 33198 42044
rect 305730 42032 305736 42044
rect 305788 42032 305794 42084
rect 38654 40740 38660 40792
rect 38712 40780 38718 40792
rect 280890 40780 280896 40792
rect 38712 40752 280896 40780
rect 38712 40740 38718 40752
rect 280890 40740 280896 40752
rect 280948 40740 280954 40792
rect 11054 40672 11060 40724
rect 11112 40712 11118 40724
rect 296162 40712 296168 40724
rect 11112 40684 296168 40712
rect 11112 40672 11118 40684
rect 296162 40672 296168 40684
rect 296220 40672 296226 40724
rect 51074 39380 51080 39432
rect 51132 39420 51138 39432
rect 279510 39420 279516 39432
rect 51132 39392 279516 39420
rect 51132 39380 51138 39392
rect 279510 39380 279516 39392
rect 279568 39380 279574 39432
rect 23474 39312 23480 39364
rect 23532 39352 23538 39364
rect 283650 39352 283656 39364
rect 23532 39324 283656 39352
rect 23532 39312 23538 39324
rect 283650 39312 283656 39324
rect 283708 39312 283714 39364
rect 45554 37952 45560 38004
rect 45612 37992 45618 38004
rect 275278 37992 275284 38004
rect 45612 37964 275284 37992
rect 45612 37952 45618 37964
rect 275278 37952 275284 37964
rect 275336 37952 275342 38004
rect 6914 37884 6920 37936
rect 6972 37924 6978 37936
rect 286594 37924 286600 37936
rect 6972 37896 286600 37924
rect 6972 37884 6978 37896
rect 286594 37884 286600 37896
rect 286652 37884 286658 37936
rect 11146 36524 11152 36576
rect 11204 36564 11210 36576
rect 278222 36564 278228 36576
rect 11204 36536 278228 36564
rect 11204 36524 11210 36536
rect 278222 36524 278228 36536
rect 278280 36524 278286 36576
rect 57882 35844 57888 35896
rect 57940 35884 57946 35896
rect 251174 35884 251180 35896
rect 57940 35856 251180 35884
rect 57940 35844 57946 35856
rect 251174 35844 251180 35856
rect 251232 35844 251238 35896
rect 109034 35232 109040 35284
rect 109092 35272 109098 35284
rect 287882 35272 287888 35284
rect 109092 35244 287888 35272
rect 109092 35232 109098 35244
rect 287882 35232 287888 35244
rect 287940 35232 287946 35284
rect 4798 35164 4804 35216
rect 4856 35204 4862 35216
rect 57882 35204 57888 35216
rect 4856 35176 57888 35204
rect 4856 35164 4862 35176
rect 57882 35164 57888 35176
rect 57940 35164 57946 35216
rect 85666 35164 85672 35216
rect 85724 35204 85730 35216
rect 308582 35204 308588 35216
rect 85724 35176 308588 35204
rect 85724 35164 85730 35176
rect 308582 35164 308588 35176
rect 308640 35164 308646 35216
rect 1302 34416 1308 34468
rect 1360 34456 1366 34468
rect 249150 34456 249156 34468
rect 1360 34428 249156 34456
rect 1360 34416 1366 34428
rect 249150 34416 249156 34428
rect 249208 34416 249214 34468
rect 63494 33736 63500 33788
rect 63552 33776 63558 33788
rect 283558 33776 283564 33788
rect 63552 33748 283564 33776
rect 63552 33736 63558 33748
rect 283558 33736 283564 33748
rect 283616 33736 283622 33788
rect 14 33124 20 33176
rect 72 33164 78 33176
rect 1302 33164 1308 33176
rect 72 33136 1308 33164
rect 72 33124 78 33136
rect 1302 33124 1308 33136
rect 1360 33124 1366 33176
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 43438 33096 43444 33108
rect 3568 33068 43444 33096
rect 3568 33056 3574 33068
rect 43438 33056 43444 33068
rect 43496 33056 43502 33108
rect 77294 32444 77300 32496
rect 77352 32484 77358 32496
rect 296070 32484 296076 32496
rect 77352 32456 296076 32484
rect 77352 32444 77358 32456
rect 296070 32444 296076 32456
rect 296128 32444 296134 32496
rect 37182 32376 37188 32428
rect 37240 32416 37246 32428
rect 270494 32416 270500 32428
rect 37240 32388 270500 32416
rect 37240 32376 37246 32388
rect 270494 32376 270500 32388
rect 270552 32376 270558 32428
rect 70394 31016 70400 31068
rect 70452 31056 70458 31068
rect 287790 31056 287796 31068
rect 70452 31028 287796 31056
rect 70452 31016 70458 31028
rect 287790 31016 287796 31028
rect 287848 31016 287854 31068
rect 195238 29724 195244 29776
rect 195296 29764 195302 29776
rect 251174 29764 251180 29776
rect 195296 29736 251180 29764
rect 195296 29724 195302 29736
rect 251174 29724 251180 29736
rect 251232 29724 251238 29776
rect 2866 29656 2872 29708
rect 2924 29696 2930 29708
rect 253198 29696 253204 29708
rect 2924 29668 253204 29696
rect 2924 29656 2930 29668
rect 253198 29656 253204 29668
rect 253256 29656 253262 29708
rect 43438 29588 43444 29640
rect 43496 29628 43502 29640
rect 307110 29628 307116 29640
rect 43496 29600 307116 29628
rect 43496 29588 43502 29600
rect 307110 29588 307116 29600
rect 307168 29588 307174 29640
rect 182818 28296 182824 28348
rect 182876 28336 182882 28348
rect 262214 28336 262220 28348
rect 182876 28308 262220 28336
rect 182876 28296 182882 28308
rect 262214 28296 262220 28308
rect 262272 28296 262278 28348
rect 8294 28228 8300 28280
rect 8352 28268 8358 28280
rect 301498 28268 301504 28280
rect 8352 28240 301504 28268
rect 8352 28228 8358 28240
rect 301498 28228 301504 28240
rect 301556 28228 301562 28280
rect 118694 26936 118700 26988
rect 118752 26976 118758 26988
rect 297450 26976 297456 26988
rect 118752 26948 297456 26976
rect 118752 26936 118758 26948
rect 297450 26936 297456 26948
rect 297508 26936 297514 26988
rect 59354 26868 59360 26920
rect 59412 26908 59418 26920
rect 265618 26908 265624 26920
rect 59412 26880 265624 26908
rect 59412 26868 59418 26880
rect 265618 26868 265624 26880
rect 265676 26868 265682 26920
rect 120074 25644 120080 25696
rect 120132 25684 120138 25696
rect 250438 25684 250444 25696
rect 120132 25656 250444 25684
rect 120132 25644 120138 25656
rect 250438 25644 250444 25656
rect 250496 25644 250502 25696
rect 86954 25576 86960 25628
rect 87012 25616 87018 25628
rect 297358 25616 297364 25628
rect 87012 25588 297364 25616
rect 87012 25576 87018 25588
rect 297358 25576 297364 25588
rect 297416 25576 297422 25628
rect 57974 25508 57980 25560
rect 58032 25548 58038 25560
rect 304350 25548 304356 25560
rect 58032 25520 304356 25548
rect 58032 25508 58038 25520
rect 304350 25508 304356 25520
rect 304408 25508 304414 25560
rect 204990 24216 204996 24268
rect 205048 24256 205054 24268
rect 244274 24256 244280 24268
rect 205048 24228 244280 24256
rect 205048 24216 205054 24228
rect 244274 24216 244280 24228
rect 244332 24216 244338 24268
rect 193858 24148 193864 24200
rect 193916 24188 193922 24200
rect 292574 24188 292580 24200
rect 193916 24160 292580 24188
rect 193916 24148 193922 24160
rect 292574 24148 292580 24160
rect 292632 24148 292638 24200
rect 102134 24080 102140 24132
rect 102192 24120 102198 24132
rect 272518 24120 272524 24132
rect 102192 24092 272524 24120
rect 102192 24080 102198 24092
rect 272518 24080 272524 24092
rect 272576 24080 272582 24132
rect 69106 22788 69112 22840
rect 69164 22828 69170 22840
rect 291838 22828 291844 22840
rect 69164 22800 291844 22828
rect 69164 22788 69170 22800
rect 291838 22788 291844 22800
rect 291896 22788 291902 22840
rect 19334 22720 19340 22772
rect 19392 22760 19398 22772
rect 261478 22760 261484 22772
rect 19392 22732 261484 22760
rect 19392 22720 19398 22732
rect 261478 22720 261484 22732
rect 261536 22720 261542 22772
rect 189718 21496 189724 21548
rect 189776 21536 189782 21548
rect 309134 21536 309140 21548
rect 189776 21508 309140 21536
rect 189776 21496 189782 21508
rect 309134 21496 309140 21508
rect 309192 21496 309198 21548
rect 62114 21428 62120 21480
rect 62172 21468 62178 21480
rect 300118 21468 300124 21480
rect 62172 21440 300124 21468
rect 62172 21428 62178 21440
rect 300118 21428 300124 21440
rect 300176 21428 300182 21480
rect 34422 21360 34428 21412
rect 34480 21400 34486 21412
rect 280154 21400 280160 21412
rect 34480 21372 280160 21400
rect 34480 21360 34486 21372
rect 280154 21360 280160 21372
rect 280212 21360 280218 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 40678 20652 40684 20664
rect 3476 20624 40684 20652
rect 3476 20612 3482 20624
rect 40678 20612 40684 20624
rect 40736 20612 40742 20664
rect 91094 19932 91100 19984
rect 91152 19972 91158 19984
rect 266998 19972 267004 19984
rect 91152 19944 267004 19972
rect 91152 19932 91158 19944
rect 266998 19932 267004 19944
rect 267056 19932 267062 19984
rect 191098 18708 191104 18760
rect 191156 18748 191162 18760
rect 241514 18748 241520 18760
rect 191156 18720 241520 18748
rect 191156 18708 191162 18720
rect 241514 18708 241520 18720
rect 241572 18708 241578 18760
rect 35986 18640 35992 18692
rect 36044 18680 36050 18692
rect 267090 18680 267096 18692
rect 36044 18652 267096 18680
rect 36044 18640 36050 18652
rect 267090 18640 267096 18652
rect 267148 18640 267154 18692
rect 55214 18572 55220 18624
rect 55272 18612 55278 18624
rect 298830 18612 298836 18624
rect 55272 18584 298836 18612
rect 55272 18572 55278 18584
rect 298830 18572 298836 18584
rect 298888 18572 298894 18624
rect 64782 17348 64788 17400
rect 64840 17388 64846 17400
rect 242986 17388 242992 17400
rect 64840 17360 242992 17388
rect 64840 17348 64846 17360
rect 242986 17348 242992 17360
rect 243044 17348 243050 17400
rect 111794 17280 111800 17332
rect 111852 17320 111858 17332
rect 302878 17320 302884 17332
rect 111852 17292 302884 17320
rect 111852 17280 111858 17292
rect 302878 17280 302884 17292
rect 302936 17280 302942 17332
rect 74534 17212 74540 17264
rect 74592 17252 74598 17264
rect 295978 17252 295984 17264
rect 74592 17224 295984 17252
rect 74592 17212 74598 17224
rect 295978 17212 295984 17224
rect 296036 17212 296042 17264
rect 195422 15988 195428 16040
rect 195480 16028 195486 16040
rect 295610 16028 295616 16040
rect 195480 16000 295616 16028
rect 195480 15988 195486 16000
rect 295610 15988 295616 16000
rect 295668 15988 295674 16040
rect 209130 15920 209136 15972
rect 209188 15960 209194 15972
rect 322934 15960 322940 15972
rect 209188 15932 322940 15960
rect 209188 15920 209194 15932
rect 322934 15920 322940 15932
rect 322992 15920 322998 15972
rect 48498 15852 48504 15904
rect 48556 15892 48562 15904
rect 268378 15892 268384 15904
rect 48556 15864 268384 15892
rect 48556 15852 48562 15864
rect 268378 15852 268384 15864
rect 268436 15852 268442 15904
rect 192478 14560 192484 14612
rect 192536 14600 192542 14612
rect 306374 14600 306380 14612
rect 192536 14572 306380 14600
rect 192536 14560 192542 14572
rect 306374 14560 306380 14572
rect 306432 14560 306438 14612
rect 40218 14492 40224 14544
rect 40276 14532 40282 14544
rect 257338 14532 257344 14544
rect 40276 14504 257344 14532
rect 40276 14492 40282 14504
rect 257338 14492 257344 14504
rect 257396 14492 257402 14544
rect 54938 14424 54944 14476
rect 54996 14464 55002 14476
rect 290458 14464 290464 14476
rect 54996 14436 290464 14464
rect 54996 14424 55002 14436
rect 290458 14424 290464 14436
rect 290516 14424 290522 14476
rect 216214 13132 216220 13184
rect 216272 13172 216278 13184
rect 259454 13172 259460 13184
rect 216272 13144 259460 13172
rect 216272 13132 216278 13144
rect 259454 13132 259460 13144
rect 259512 13132 259518 13184
rect 203518 13064 203524 13116
rect 203576 13104 203582 13116
rect 267734 13104 267740 13116
rect 203576 13076 267740 13104
rect 203576 13064 203582 13076
rect 267734 13064 267740 13076
rect 267792 13064 267798 13116
rect 187050 11840 187056 11892
rect 187108 11880 187114 11892
rect 247586 11880 247592 11892
rect 187108 11852 247592 11880
rect 187108 11840 187114 11852
rect 247586 11840 247592 11852
rect 247644 11840 247650 11892
rect 191190 11772 191196 11824
rect 191248 11812 191254 11824
rect 327994 11812 328000 11824
rect 191248 11784 328000 11812
rect 191248 11772 191254 11784
rect 327994 11772 328000 11784
rect 328052 11772 328058 11824
rect 80882 11704 80888 11756
rect 80940 11744 80946 11756
rect 286410 11744 286416 11756
rect 80940 11716 286416 11744
rect 80940 11704 80946 11716
rect 286410 11704 286416 11716
rect 286468 11704 286474 11756
rect 186958 10412 186964 10464
rect 187016 10452 187022 10464
rect 256694 10452 256700 10464
rect 187016 10424 256700 10452
rect 187016 10412 187022 10424
rect 256694 10412 256700 10424
rect 256752 10412 256758 10464
rect 52546 10344 52552 10396
rect 52604 10384 52610 10396
rect 264238 10384 264244 10396
rect 52604 10356 264244 10384
rect 52604 10344 52610 10356
rect 264238 10344 264244 10356
rect 264296 10344 264302 10396
rect 44266 10276 44272 10328
rect 44324 10316 44330 10328
rect 289170 10316 289176 10328
rect 44324 10288 289176 10316
rect 44324 10276 44330 10288
rect 289170 10276 289176 10288
rect 289228 10276 289234 10328
rect 200758 9052 200764 9104
rect 200816 9092 200822 9104
rect 254670 9092 254676 9104
rect 200816 9064 254676 9092
rect 200816 9052 200822 9064
rect 254670 9052 254676 9064
rect 254728 9052 254734 9104
rect 119890 8984 119896 9036
rect 119948 9024 119954 9036
rect 298738 9024 298744 9036
rect 119948 8996 298744 9024
rect 119948 8984 119954 8996
rect 298738 8984 298744 8996
rect 298796 8984 298802 9036
rect 41874 8916 41880 8968
rect 41932 8956 41938 8968
rect 307018 8956 307024 8968
rect 41932 8928 307024 8956
rect 41932 8916 41938 8928
rect 307018 8916 307024 8928
rect 307076 8916 307082 8968
rect 216030 7692 216036 7744
rect 216088 7732 216094 7744
rect 239306 7732 239312 7744
rect 216088 7704 239312 7732
rect 216088 7692 216094 7704
rect 239306 7692 239312 7704
rect 239364 7692 239370 7744
rect 39942 7624 39948 7676
rect 40000 7664 40006 7676
rect 168374 7664 168380 7676
rect 40000 7636 168380 7664
rect 40000 7624 40006 7636
rect 168374 7624 168380 7636
rect 168432 7624 168438 7676
rect 197998 7624 198004 7676
rect 198056 7664 198062 7676
rect 249978 7664 249984 7676
rect 198056 7636 249984 7664
rect 198056 7624 198062 7636
rect 249978 7624 249984 7636
rect 250036 7624 250042 7676
rect 4062 7556 4068 7608
rect 4120 7596 4126 7608
rect 25498 7596 25504 7608
rect 4120 7568 25504 7596
rect 4120 7556 4126 7568
rect 25498 7556 25504 7568
rect 25556 7556 25562 7608
rect 105722 7556 105728 7608
rect 105780 7596 105786 7608
rect 289078 7596 289084 7608
rect 105780 7568 289084 7596
rect 105780 7556 105786 7568
rect 289078 7556 289084 7568
rect 289136 7556 289142 7608
rect 199378 6264 199384 6316
rect 199436 6304 199442 6316
rect 292574 6304 292580 6316
rect 199436 6276 292580 6304
rect 199436 6264 199442 6276
rect 292574 6264 292580 6276
rect 292632 6264 292638 6316
rect 65518 6196 65524 6248
rect 65576 6236 65582 6248
rect 305638 6236 305644 6248
rect 65576 6208 305644 6236
rect 65576 6196 65582 6208
rect 305638 6196 305644 6208
rect 305696 6196 305702 6248
rect 19426 6128 19432 6180
rect 19484 6168 19490 6180
rect 282178 6168 282184 6180
rect 19484 6140 282184 6168
rect 19484 6128 19490 6140
rect 282178 6128 282184 6140
rect 282236 6128 282242 6180
rect 117590 4836 117596 4888
rect 117648 4876 117654 4888
rect 278130 4876 278136 4888
rect 117648 4848 278136 4876
rect 117648 4836 117654 4848
rect 278130 4836 278136 4848
rect 278188 4836 278194 4888
rect 62022 4768 62028 4820
rect 62080 4808 62086 4820
rect 258718 4808 258724 4820
rect 62080 4780 258724 4808
rect 62080 4768 62086 4780
rect 258718 4768 258724 4780
rect 258776 4768 258782 4820
rect 309686 4088 309692 4140
rect 309744 4128 309750 4140
rect 318518 4128 318524 4140
rect 309744 4100 318524 4128
rect 309744 4088 309750 4100
rect 318518 4088 318524 4100
rect 318576 4088 318582 4140
rect 320910 3720 320916 3732
rect 316006 3692 320916 3720
rect 217318 3612 217324 3664
rect 217376 3652 217382 3664
rect 242894 3652 242900 3664
rect 217376 3624 242900 3652
rect 217376 3612 217382 3624
rect 242894 3612 242900 3624
rect 242952 3612 242958 3664
rect 308398 3612 308404 3664
rect 308456 3652 308462 3664
rect 316006 3652 316034 3692
rect 320910 3680 320916 3692
rect 320968 3680 320974 3732
rect 308456 3624 316034 3652
rect 308456 3612 308462 3624
rect 316126 3612 316132 3664
rect 316184 3652 316190 3664
rect 317322 3652 317328 3664
rect 316184 3624 317328 3652
rect 316184 3612 316190 3624
rect 317322 3612 317328 3624
rect 317380 3612 317386 3664
rect 1670 3544 1676 3596
rect 1728 3584 1734 3596
rect 4798 3584 4804 3596
rect 1728 3556 4804 3584
rect 1728 3544 1734 3556
rect 4798 3544 4804 3556
rect 4856 3544 4862 3596
rect 125870 3544 125876 3596
rect 125928 3584 125934 3596
rect 171134 3584 171140 3596
rect 125928 3556 171140 3584
rect 125928 3544 125934 3556
rect 171134 3544 171140 3556
rect 171192 3544 171198 3596
rect 213178 3544 213184 3596
rect 213236 3584 213242 3596
rect 240502 3584 240508 3596
rect 213236 3556 240508 3584
rect 213236 3544 213242 3556
rect 240502 3544 240508 3556
rect 240560 3544 240566 3596
rect 251174 3544 251180 3596
rect 251232 3584 251238 3596
rect 252370 3584 252376 3596
rect 251232 3556 252376 3584
rect 251232 3544 251238 3556
rect 252370 3544 252376 3556
rect 252428 3544 252434 3596
rect 259454 3544 259460 3596
rect 259512 3584 259518 3596
rect 260650 3584 260656 3596
rect 259512 3556 260656 3584
rect 259512 3544 259518 3556
rect 260650 3544 260656 3556
rect 260708 3544 260714 3596
rect 299474 3544 299480 3596
rect 299532 3584 299538 3596
rect 300762 3584 300768 3596
rect 299532 3556 300768 3584
rect 299532 3544 299538 3556
rect 300762 3544 300768 3556
rect 300820 3544 300826 3596
rect 307846 3544 307852 3596
rect 307904 3584 307910 3596
rect 309042 3584 309048 3596
rect 307904 3556 309048 3584
rect 307904 3544 307910 3556
rect 309042 3544 309048 3556
rect 309100 3544 309106 3596
rect 309870 3544 309876 3596
rect 309928 3584 309934 3596
rect 329190 3584 329196 3596
rect 309928 3556 329196 3584
rect 309928 3544 309934 3556
rect 329190 3544 329196 3556
rect 329248 3544 329254 3596
rect 11054 3476 11060 3528
rect 11112 3516 11118 3528
rect 11974 3516 11980 3528
rect 11112 3488 11980 3516
rect 11112 3476 11118 3488
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 25314 3476 25320 3528
rect 25372 3516 25378 3528
rect 43438 3516 43444 3528
rect 25372 3488 43444 3516
rect 25372 3476 25378 3488
rect 43438 3476 43444 3488
rect 43496 3476 43502 3528
rect 44174 3476 44180 3528
rect 44232 3516 44238 3528
rect 45094 3516 45100 3528
rect 44232 3488 45100 3516
rect 44232 3476 44238 3488
rect 45094 3476 45100 3488
rect 45152 3476 45158 3528
rect 52454 3476 52460 3528
rect 52512 3516 52518 3528
rect 53374 3516 53380 3528
rect 52512 3488 53380 3516
rect 52512 3476 52518 3488
rect 53374 3476 53380 3488
rect 53432 3476 53438 3528
rect 85574 3476 85580 3528
rect 85632 3516 85638 3528
rect 86494 3516 86500 3528
rect 85632 3488 86500 3516
rect 85632 3476 85638 3488
rect 86494 3476 86500 3488
rect 86552 3476 86558 3528
rect 103330 3476 103336 3528
rect 103388 3516 103394 3528
rect 188338 3516 188344 3528
rect 103388 3488 188344 3516
rect 103388 3476 103394 3488
rect 188338 3476 188344 3488
rect 188396 3476 188402 3528
rect 215938 3476 215944 3528
rect 215996 3516 216002 3528
rect 253474 3516 253480 3528
rect 215996 3488 253480 3516
rect 215996 3476 216002 3488
rect 253474 3476 253480 3488
rect 253532 3476 253538 3528
rect 287698 3476 287704 3528
rect 287756 3516 287762 3528
rect 312630 3516 312636 3528
rect 287756 3488 312636 3516
rect 287756 3476 287762 3488
rect 312630 3476 312636 3488
rect 312688 3476 312694 3528
rect 324406 3476 324412 3528
rect 324464 3516 324470 3528
rect 325602 3516 325608 3528
rect 324464 3488 325608 3516
rect 324464 3476 324470 3488
rect 325602 3476 325608 3488
rect 325660 3476 325666 3528
rect 349154 3476 349160 3528
rect 349212 3516 349218 3528
rect 350442 3516 350448 3528
rect 349212 3488 350448 3516
rect 349212 3476 349218 3488
rect 350442 3476 350448 3488
rect 350500 3476 350506 3528
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 15194 3448 15200 3460
rect 6512 3420 15200 3448
rect 6512 3408 6518 3420
rect 15194 3408 15200 3420
rect 15252 3408 15258 3460
rect 43070 3408 43076 3460
rect 43128 3448 43134 3460
rect 178678 3448 178684 3460
rect 43128 3420 178684 3448
rect 43128 3408 43134 3420
rect 178678 3408 178684 3420
rect 178736 3408 178742 3460
rect 204898 3408 204904 3460
rect 204956 3448 204962 3460
rect 246390 3448 246396 3460
rect 204956 3420 246396 3448
rect 204956 3408 204962 3420
rect 246390 3408 246396 3420
rect 246448 3408 246454 3460
rect 279418 3408 279424 3460
rect 279476 3448 279482 3460
rect 311434 3448 311440 3460
rect 279476 3420 311440 3448
rect 279476 3408 279482 3420
rect 311434 3408 311440 3420
rect 311492 3408 311498 3460
rect 342162 3408 342168 3460
rect 342220 3448 342226 3460
rect 353294 3448 353300 3460
rect 342220 3420 353300 3448
rect 342220 3408 342226 3420
rect 353294 3408 353300 3420
rect 353352 3408 353358 3460
rect 235810 2932 235816 2984
rect 235868 2972 235874 2984
rect 238018 2972 238024 2984
rect 235868 2944 238024 2972
rect 235868 2932 235874 2944
rect 238018 2932 238024 2944
rect 238076 2932 238082 2984
rect 66714 2116 66720 2168
rect 66772 2156 66778 2168
rect 304258 2156 304264 2168
rect 66772 2128 304264 2156
rect 66772 2116 66778 2128
rect 304258 2116 304264 2128
rect 304316 2116 304322 2168
rect 15930 2048 15936 2100
rect 15988 2088 15994 2100
rect 291930 2088 291936 2100
rect 15988 2060 291936 2088
rect 15988 2048 15994 2060
rect 291930 2048 291936 2060
rect 291988 2048 291994 2100
<< via1 >>
rect 201500 703128 201552 703180
rect 202788 703128 202840 703180
rect 98644 703060 98696 703112
rect 332508 703060 332560 703112
rect 79324 702992 79376 703044
rect 364984 702992 365036 703044
rect 106280 702924 106332 702976
rect 413652 702924 413704 702976
rect 117228 702856 117280 702908
rect 462320 702856 462372 702908
rect 79416 702788 79468 702840
rect 429844 702788 429896 702840
rect 123484 702720 123536 702772
rect 478512 702720 478564 702772
rect 119988 702652 120040 702704
rect 494796 702652 494848 702704
rect 115848 702584 115900 702636
rect 559656 702584 559708 702636
rect 81348 702516 81400 702568
rect 527180 702516 527232 702568
rect 57244 702448 57296 702500
rect 543464 702448 543516 702500
rect 86224 700340 86276 700392
rect 154120 700340 154172 700392
rect 155224 700340 155276 700392
rect 218980 700340 219032 700392
rect 66168 700272 66220 700324
rect 170312 700272 170364 700324
rect 220084 700272 220136 700324
rect 235172 700272 235224 700324
rect 341524 700272 341576 700324
rect 348792 700272 348844 700324
rect 8116 700204 8168 700256
rect 14464 700204 14516 700256
rect 395344 699660 395396 699712
rect 397460 699660 397512 699712
rect 24308 698912 24360 698964
rect 110420 698912 110472 698964
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 68284 694764 68336 694816
rect 282920 694764 282972 694816
rect 3424 683136 3476 683188
rect 75184 683136 75236 683188
rect 3516 670692 3568 670744
rect 58624 670692 58676 670744
rect 87604 670692 87656 670744
rect 580172 670692 580224 670744
rect 3424 656888 3476 656940
rect 35164 656888 35216 656940
rect 142804 643084 142856 643136
rect 580172 643084 580224 643136
rect 124864 630640 124916 630692
rect 579988 630640 580040 630692
rect 3516 618264 3568 618316
rect 15844 618264 15896 618316
rect 3516 605820 3568 605872
rect 25504 605820 25556 605872
rect 146944 590656 146996 590708
rect 580172 590656 580224 590708
rect 3332 579640 3384 579692
rect 32404 579640 32456 579692
rect 70308 576852 70360 576904
rect 580172 576852 580224 576904
rect 3240 565836 3292 565888
rect 60740 565836 60792 565888
rect 148324 563048 148376 563100
rect 580172 563048 580224 563100
rect 3516 553800 3568 553852
rect 7564 553800 7616 553852
rect 122104 536800 122156 536852
rect 579896 536800 579948 536852
rect 7564 530544 7616 530596
rect 111800 530544 111852 530596
rect 2964 527144 3016 527196
rect 7564 527144 7616 527196
rect 141424 524424 141476 524476
rect 580172 524424 580224 524476
rect 3516 514768 3568 514820
rect 101404 514768 101456 514820
rect 76564 510620 76616 510672
rect 580172 510620 580224 510672
rect 3056 500964 3108 501016
rect 93124 500964 93176 501016
rect 126244 484372 126296 484424
rect 580172 484372 580224 484424
rect 3056 474716 3108 474768
rect 35256 474716 35308 474768
rect 116584 470568 116636 470620
rect 580172 470568 580224 470620
rect 2780 462544 2832 462596
rect 4804 462544 4856 462596
rect 97264 456764 97316 456816
rect 580172 456764 580224 456816
rect 35164 453296 35216 453348
rect 90364 453296 90416 453348
rect 3148 448536 3200 448588
rect 11704 448536 11756 448588
rect 130384 430584 130436 430636
rect 579896 430584 579948 430636
rect 3516 422288 3568 422340
rect 108304 422288 108356 422340
rect 72424 418140 72476 418192
rect 580172 418140 580224 418192
rect 2872 409844 2924 409896
rect 110604 409844 110656 409896
rect 97356 404336 97408 404388
rect 580172 404336 580224 404388
rect 68836 403588 68888 403640
rect 220084 403588 220136 403640
rect 15844 400868 15896 400920
rect 42800 400868 42852 400920
rect 42800 400188 42852 400240
rect 44088 400188 44140 400240
rect 99380 400188 99432 400240
rect 14464 399440 14516 399492
rect 40868 399440 40920 399492
rect 91744 399440 91796 399492
rect 97264 399440 97316 399492
rect 40868 398828 40920 398880
rect 41328 398828 41380 398880
rect 89720 398828 89772 398880
rect 68744 398080 68796 398132
rect 86224 398080 86276 398132
rect 3516 397468 3568 397520
rect 15200 397468 15252 397520
rect 15200 396720 15252 396772
rect 48228 396720 48280 396772
rect 48228 396040 48280 396092
rect 111984 396040 112036 396092
rect 71044 395292 71096 395344
rect 136640 395292 136692 395344
rect 135260 393932 135312 393984
rect 266360 393932 266412 393984
rect 81532 393320 81584 393372
rect 135260 393320 135312 393372
rect 115204 392572 115256 392624
rect 299480 392572 299532 392624
rect 7564 391212 7616 391264
rect 111892 391212 111944 391264
rect 118608 391212 118660 391264
rect 201500 391212 201552 391264
rect 75000 390532 75052 390584
rect 166264 390532 166316 390584
rect 112444 389784 112496 389836
rect 148324 389784 148376 389836
rect 108304 389308 108356 389360
rect 109684 389308 109736 389360
rect 65984 389240 66036 389292
rect 232504 389240 232556 389292
rect 70400 389172 70452 389224
rect 353300 389172 353352 389224
rect 88340 388424 88392 388476
rect 117320 388424 117372 388476
rect 137100 388424 137152 388476
rect 155224 388424 155276 388476
rect 102140 387880 102192 387932
rect 136824 387880 136876 387932
rect 137100 387880 137152 387932
rect 85672 387812 85724 387864
rect 169024 387812 169076 387864
rect 104900 387744 104952 387796
rect 110696 387744 110748 387796
rect 40040 387064 40092 387116
rect 51080 387064 51132 387116
rect 76656 387064 76708 387116
rect 97356 387064 97408 387116
rect 113916 387064 113968 387116
rect 580264 387064 580316 387116
rect 51080 386520 51132 386572
rect 52368 386520 52420 386572
rect 76748 386520 76800 386572
rect 100760 386520 100812 386572
rect 101404 386520 101456 386572
rect 147680 386520 147732 386572
rect 68836 386452 68888 386504
rect 132500 386452 132552 386504
rect 73712 386384 73764 386436
rect 313924 386384 313976 386436
rect 84936 386316 84988 386368
rect 87604 386316 87656 386368
rect 109684 385364 109736 385416
rect 124220 385364 124272 385416
rect 88248 385296 88300 385348
rect 121460 385296 121512 385348
rect 90364 385228 90416 385280
rect 125600 385228 125652 385280
rect 81348 385160 81400 385212
rect 128544 385160 128596 385212
rect 57796 385092 57848 385144
rect 98644 385092 98696 385144
rect 100668 385092 100720 385144
rect 160744 385092 160796 385144
rect 70216 385024 70268 385076
rect 76564 385024 76616 385076
rect 94596 385024 94648 385076
rect 309784 385024 309836 385076
rect 68376 384140 68428 384192
rect 72424 384140 72476 384192
rect 96528 383936 96580 383988
rect 128360 383936 128412 383988
rect 93124 383868 93176 383920
rect 132592 383868 132644 383920
rect 73068 383800 73120 383852
rect 118700 383800 118752 383852
rect 49608 383732 49660 383784
rect 71044 383732 71096 383784
rect 97908 383732 97960 383784
rect 195244 383732 195296 383784
rect 62028 383664 62080 383716
rect 84936 383664 84988 383716
rect 103888 383664 103940 383716
rect 215944 383664 215996 383716
rect 84568 382916 84620 382968
rect 100668 382916 100720 382968
rect 101864 382644 101916 382696
rect 209044 382644 209096 382696
rect 77852 382576 77904 382628
rect 79416 382576 79468 382628
rect 96160 382576 96212 382628
rect 280804 382576 280856 382628
rect 59268 382508 59320 382560
rect 70216 382508 70268 382560
rect 60648 382440 60700 382492
rect 76656 382508 76708 382560
rect 87696 382508 87748 382560
rect 109868 382508 109920 382560
rect 55128 382372 55180 382424
rect 77852 382440 77904 382492
rect 80704 382440 80756 382492
rect 106832 382440 106884 382492
rect 74816 382372 74868 382424
rect 89812 382372 89864 382424
rect 92848 382372 92900 382424
rect 133972 382372 134024 382424
rect 56416 382304 56468 382356
rect 81900 382304 81952 382356
rect 85304 382304 85356 382356
rect 104808 382304 104860 382356
rect 21364 382236 21416 382288
rect 72056 382236 72108 382288
rect 73068 382236 73120 382288
rect 106188 382236 106240 382288
rect 113824 382236 113876 382288
rect 74908 382168 74960 382220
rect 75184 382168 75236 382220
rect 97448 381080 97500 381132
rect 109776 381080 109828 381132
rect 50988 381012 51040 381064
rect 79324 381012 79376 381064
rect 104624 381012 104676 381064
rect 136640 381012 136692 381064
rect 74908 380944 74960 380996
rect 122840 380944 122892 380996
rect 50896 380876 50948 380928
rect 111800 380876 111852 380928
rect 112168 380876 112220 380928
rect 106832 380196 106884 380248
rect 131212 380196 131264 380248
rect 104808 380128 104860 380180
rect 173164 380128 173216 380180
rect 66076 380060 66128 380112
rect 71964 380060 72016 380112
rect 71688 379720 71740 379772
rect 109500 379720 109552 379772
rect 34336 379652 34388 379704
rect 78772 379652 78824 379704
rect 53656 379584 53708 379636
rect 99932 379584 99984 379636
rect 103152 379584 103204 379636
rect 121552 379584 121604 379636
rect 43996 379516 44048 379568
rect 105084 379516 105136 379568
rect 107016 379516 107068 379568
rect 114652 379516 114704 379568
rect 107660 379448 107712 379500
rect 109684 379448 109736 379500
rect 71688 379380 71740 379432
rect 73712 379380 73764 379432
rect 108304 379244 108356 379296
rect 111800 378428 111852 378480
rect 114008 378428 114060 378480
rect 140780 378156 140832 378208
rect 39948 376796 40000 376848
rect 67640 376796 67692 376848
rect 111800 376796 111852 376848
rect 119344 376796 119396 376848
rect 35808 376728 35860 376780
rect 67732 376728 67784 376780
rect 115756 376728 115808 376780
rect 128452 376728 128504 376780
rect 111800 375708 111852 375760
rect 115756 375708 115808 375760
rect 64788 375368 64840 375420
rect 67640 375368 67692 375420
rect 112076 375368 112128 375420
rect 116676 375368 116728 375420
rect 3516 374620 3568 374672
rect 67548 374620 67600 374672
rect 53748 374008 53800 374060
rect 57244 374008 57296 374060
rect 111800 374008 111852 374060
rect 196624 374008 196676 374060
rect 67640 373940 67692 373992
rect 114008 373260 114060 373312
rect 349160 373260 349212 373312
rect 111984 372784 112036 372836
rect 112168 372784 112220 372836
rect 65984 372512 66036 372564
rect 67640 372512 67692 372564
rect 112352 372512 112404 372564
rect 113916 372512 113968 372564
rect 3332 371220 3384 371272
rect 39304 371220 39356 371272
rect 67272 371220 67324 371272
rect 68652 371220 68704 371272
rect 109684 370472 109736 370524
rect 271880 370472 271932 370524
rect 111800 369928 111852 369980
rect 114468 369928 114520 369980
rect 112352 369112 112404 369164
rect 120080 369112 120132 369164
rect 60464 368500 60516 368552
rect 67640 368500 67692 368552
rect 37188 367072 37240 367124
rect 67640 367072 67692 367124
rect 111800 367072 111852 367124
rect 324964 367072 325016 367124
rect 63408 365712 63460 365764
rect 67640 365712 67692 365764
rect 109316 365712 109368 365764
rect 110328 365712 110380 365764
rect 118608 365712 118660 365764
rect 111800 364760 111852 364812
rect 114560 364760 114612 364812
rect 111800 364624 111852 364676
rect 112076 364624 112128 364676
rect 63316 364420 63368 364472
rect 67640 364420 67692 364472
rect 59176 364352 59228 364404
rect 67732 364352 67784 364404
rect 111984 364352 112036 364404
rect 142160 364352 142212 364404
rect 316776 364352 316828 364404
rect 579620 364352 579672 364404
rect 119344 363604 119396 363656
rect 282920 363604 282972 363656
rect 111892 362244 111944 362296
rect 122104 362244 122156 362296
rect 111984 362176 112036 362228
rect 116584 362176 116636 362228
rect 118608 362176 118660 362228
rect 580356 362176 580408 362228
rect 34428 361564 34480 361616
rect 67640 361564 67692 361616
rect 109592 361496 109644 361548
rect 123484 361496 123536 361548
rect 61844 360272 61896 360324
rect 67732 360272 67784 360324
rect 68284 360272 68336 360324
rect 111892 360272 111944 360324
rect 202144 360272 202196 360324
rect 48136 360204 48188 360256
rect 67640 360204 67692 360256
rect 111892 358844 111944 358896
rect 122932 358844 122984 358896
rect 37096 358776 37148 358828
rect 67640 358776 67692 358828
rect 111984 358776 112036 358828
rect 186964 358776 187016 358828
rect 57888 357484 57940 357536
rect 67732 357484 67784 357536
rect 3332 357416 3384 357468
rect 22744 357416 22796 357468
rect 56508 357416 56560 357468
rect 67640 357416 67692 357468
rect 111892 357348 111944 357400
rect 118516 357416 118568 357468
rect 127072 357416 127124 357468
rect 55036 356056 55088 356108
rect 67640 356056 67692 356108
rect 111892 356056 111944 356108
rect 211804 356056 211856 356108
rect 60556 354764 60608 354816
rect 66168 354764 66220 354816
rect 67732 354764 67784 354816
rect 64604 354696 64656 354748
rect 67640 354696 67692 354748
rect 111892 354696 111944 354748
rect 206284 354696 206336 354748
rect 65984 353336 66036 353388
rect 68100 353336 68152 353388
rect 46848 353268 46900 353320
rect 67640 353268 67692 353320
rect 111892 353268 111944 353320
rect 139400 353268 139452 353320
rect 61936 351908 61988 351960
rect 67640 351908 67692 351960
rect 111064 351908 111116 351960
rect 129740 351908 129792 351960
rect 42708 350548 42760 350600
rect 67640 350548 67692 350600
rect 111892 350548 111944 350600
rect 143540 350548 143592 350600
rect 146944 350548 146996 350600
rect 112168 349188 112220 349240
rect 135168 349188 135220 349240
rect 111892 349120 111944 349172
rect 269764 349120 269816 349172
rect 135168 348372 135220 348424
rect 346400 348372 346452 348424
rect 64696 347828 64748 347880
rect 67640 347828 67692 347880
rect 45468 347760 45520 347812
rect 67732 347760 67784 347812
rect 111892 347760 111944 347812
rect 206376 347760 206428 347812
rect 111892 346400 111944 346452
rect 278044 346400 278096 346452
rect 3332 346332 3384 346384
rect 21364 346332 21416 346384
rect 111892 345108 111944 345160
rect 123024 345108 123076 345160
rect 112168 345040 112220 345092
rect 216036 345040 216088 345092
rect 60740 344972 60792 345024
rect 67640 344972 67692 345024
rect 22744 344292 22796 344344
rect 51080 344292 51132 344344
rect 54944 344292 54996 344344
rect 60740 344292 60792 344344
rect 111984 344224 112036 344276
rect 112168 344224 112220 344276
rect 111892 343816 111944 343868
rect 115848 343816 115900 343868
rect 51080 343612 51132 343664
rect 52184 343612 52236 343664
rect 67732 343612 67784 343664
rect 111984 343612 112036 343664
rect 316684 343612 316736 343664
rect 111892 343544 111944 343596
rect 119988 343544 120040 343596
rect 115848 342864 115900 342916
rect 277400 342864 277452 342916
rect 111892 342184 111944 342236
rect 117228 342184 117280 342236
rect 124956 341504 125008 341556
rect 580264 341504 580316 341556
rect 65892 340892 65944 340944
rect 67640 340892 67692 340944
rect 117228 340892 117280 340944
rect 120724 340892 120776 340944
rect 110328 340144 110380 340196
rect 112168 340144 112220 340196
rect 70492 339940 70544 339992
rect 79324 339940 79376 339992
rect 107568 339940 107620 339992
rect 395344 340144 395396 340196
rect 4804 339396 4856 339448
rect 83556 339396 83608 339448
rect 84844 339396 84896 339448
rect 316776 339396 316828 339448
rect 65984 339328 66036 339380
rect 125692 339328 125744 339380
rect 126244 339328 126296 339380
rect 58624 339260 58676 339312
rect 91100 339260 91152 339312
rect 91928 339260 91980 339312
rect 95148 339260 95200 339312
rect 117320 339260 117372 339312
rect 106280 338852 106332 338904
rect 109592 338852 109644 338904
rect 105544 338784 105596 338836
rect 113364 338784 113416 338836
rect 68560 338716 68612 338768
rect 284300 338716 284352 338768
rect 32404 338036 32456 338088
rect 98644 338036 98696 338088
rect 104164 338036 104216 338088
rect 115204 338036 115256 338088
rect 66076 337968 66128 338020
rect 73896 337968 73948 338020
rect 78404 337968 78456 338020
rect 129832 338036 129884 338088
rect 130384 338036 130436 338088
rect 80980 337900 81032 337952
rect 107568 337900 107620 337952
rect 84200 337832 84252 337884
rect 90088 337832 90140 337884
rect 70676 337696 70728 337748
rect 72424 337696 72476 337748
rect 100300 337696 100352 337748
rect 101404 337696 101456 337748
rect 71320 337560 71372 337612
rect 73804 337560 73856 337612
rect 87420 337560 87472 337612
rect 89076 337560 89128 337612
rect 100024 337560 100076 337612
rect 114560 337560 114612 337612
rect 109316 337492 109368 337544
rect 191104 337492 191156 337544
rect 73252 337424 73304 337476
rect 80428 337424 80480 337476
rect 81624 337424 81676 337476
rect 188344 337424 188396 337476
rect 74540 337356 74592 337408
rect 87604 337356 87656 337408
rect 92572 337356 92624 337408
rect 307024 337356 307076 337408
rect 70032 336948 70084 337000
rect 75276 336948 75328 337000
rect 72608 336744 72660 336796
rect 75184 336744 75236 336796
rect 35256 336676 35308 336728
rect 95884 336676 95936 336728
rect 96436 336676 96488 336728
rect 68836 336132 68888 336184
rect 269120 336132 269172 336184
rect 60464 336064 60516 336116
rect 88984 336064 89036 336116
rect 90088 336064 90140 336116
rect 343640 336064 343692 336116
rect 88708 335996 88760 336048
rect 126980 335996 127032 336048
rect 582380 335996 582432 336048
rect 56324 334840 56376 334892
rect 82912 334840 82964 334892
rect 57704 334772 57756 334824
rect 94504 334772 94556 334824
rect 3424 334568 3476 334620
rect 53564 334568 53616 334620
rect 99656 334704 99708 334756
rect 99748 334704 99800 334756
rect 112076 334704 112128 334756
rect 131120 334704 131172 334756
rect 61936 334636 61988 334688
rect 133880 334636 133932 334688
rect 68744 334568 68796 334620
rect 309876 334568 309928 334620
rect 107384 333888 107436 333940
rect 341524 333888 341576 333940
rect 25504 333820 25556 333872
rect 107752 333820 107804 333872
rect 67364 333208 67416 333260
rect 273260 333208 273312 333260
rect 106924 332596 106976 332648
rect 107384 332596 107436 332648
rect 39304 332528 39356 332580
rect 99748 332528 99800 332580
rect 52276 331848 52328 331900
rect 91284 331848 91336 331900
rect 80428 331168 80480 331220
rect 124312 331168 124364 331220
rect 124956 331168 125008 331220
rect 61936 330556 61988 330608
rect 113272 330556 113324 330608
rect 98368 330488 98420 330540
rect 293960 330488 294012 330540
rect 67456 329196 67508 329248
rect 115204 329196 115256 329248
rect 39856 329128 39908 329180
rect 102876 329128 102928 329180
rect 69112 329060 69164 329112
rect 281540 329060 281592 329112
rect 65892 328380 65944 328432
rect 140872 328380 140924 328432
rect 141424 328380 141476 328432
rect 73160 327768 73212 327820
rect 109132 327768 109184 327820
rect 79048 327700 79100 327752
rect 204904 327700 204956 327752
rect 106740 326340 106792 326392
rect 152464 326340 152516 326392
rect 73896 324912 73948 324964
rect 114560 324912 114612 324964
rect 102140 323688 102192 323740
rect 121552 323688 121604 323740
rect 121828 323688 121880 323740
rect 97080 323620 97132 323672
rect 284392 323620 284444 323672
rect 84292 323552 84344 323604
rect 109500 323552 109552 323604
rect 121828 323552 121880 323604
rect 582564 323552 582616 323604
rect 71044 322328 71096 322380
rect 102140 322328 102192 322380
rect 93860 322260 93912 322312
rect 287060 322260 287112 322312
rect 68928 322192 68980 322244
rect 308404 322192 308456 322244
rect 101404 320832 101456 320884
rect 349252 320832 349304 320884
rect 79324 319472 79376 319524
rect 155224 319472 155276 319524
rect 59176 319404 59228 319456
rect 198004 319404 198056 319456
rect 95148 318724 95200 318776
rect 101404 318724 101456 318776
rect 77116 318044 77168 318096
rect 204996 318044 205048 318096
rect 129004 317364 129056 317416
rect 131212 317364 131264 317416
rect 580172 317364 580224 317416
rect 64604 316820 64656 316872
rect 124404 316820 124456 316872
rect 61844 316752 61896 316804
rect 134064 316752 134116 316804
rect 76472 316684 76524 316736
rect 213184 316684 213236 316736
rect 89352 315256 89404 315308
rect 146944 315256 146996 315308
rect 63132 314032 63184 314084
rect 84844 314032 84896 314084
rect 94504 313964 94556 314016
rect 108672 313964 108724 314016
rect 63408 313896 63460 313948
rect 129924 313896 129976 313948
rect 71964 312604 72016 312656
rect 287704 312604 287756 312656
rect 3424 312536 3476 312588
rect 115940 312536 115992 312588
rect 124404 312468 124456 312520
rect 124864 312468 124916 312520
rect 580172 312536 580224 312588
rect 72424 311176 72476 311228
rect 103520 311176 103572 311228
rect 79692 311108 79744 311160
rect 180064 311108 180116 311160
rect 75920 310496 75972 310548
rect 295984 310496 296036 310548
rect 75828 309816 75880 309868
rect 121644 309816 121696 309868
rect 75276 309748 75328 309800
rect 291200 309748 291252 309800
rect 101588 308660 101640 308712
rect 113824 308660 113876 308712
rect 87604 308592 87656 308644
rect 106924 308592 106976 308644
rect 89076 308524 89128 308576
rect 274640 308524 274692 308576
rect 69020 308456 69072 308508
rect 298100 308456 298152 308508
rect 80060 308388 80112 308440
rect 121460 308388 121512 308440
rect 582840 308388 582892 308440
rect 76564 307096 76616 307148
rect 159364 307096 159416 307148
rect 88064 307028 88116 307080
rect 278780 307028 278832 307080
rect 81440 306416 81492 306468
rect 246304 306416 246356 306468
rect 89720 306348 89772 306400
rect 300124 306348 300176 306400
rect 3424 306280 3476 306332
rect 42708 306280 42760 306332
rect 95884 305804 95936 305856
rect 123116 305804 123168 305856
rect 61844 305736 61896 305788
rect 110420 305736 110472 305788
rect 42708 305668 42760 305720
rect 117412 305668 117464 305720
rect 86132 305600 86184 305652
rect 217324 305600 217376 305652
rect 88340 304988 88392 305040
rect 356060 304988 356112 305040
rect 72240 304240 72292 304292
rect 124220 304240 124272 304292
rect 106096 303764 106148 303816
rect 110512 303764 110564 303816
rect 111708 303764 111760 303816
rect 111892 303764 111944 303816
rect 116676 303764 116728 303816
rect 117320 303764 117372 303816
rect 79324 303696 79376 303748
rect 229744 303696 229796 303748
rect 67456 303628 67508 303680
rect 226984 303628 227036 303680
rect 69020 302948 69072 303000
rect 111800 302948 111852 303000
rect 86776 302880 86828 302932
rect 151084 302880 151136 302932
rect 100852 302404 100904 302456
rect 244924 302404 244976 302456
rect 74540 302336 74592 302388
rect 222844 302336 222896 302388
rect 106372 302268 106424 302320
rect 319444 302268 319496 302320
rect 103612 302200 103664 302252
rect 349344 302200 349396 302252
rect 122104 302132 122156 302184
rect 124220 302132 124272 302184
rect 66076 301452 66128 301504
rect 111708 301452 111760 301504
rect 583116 301452 583168 301504
rect 102140 300976 102192 301028
rect 199384 300976 199436 301028
rect 73252 300908 73304 300960
rect 192484 300908 192536 300960
rect 85580 300840 85632 300892
rect 224224 300840 224276 300892
rect 52184 300160 52236 300212
rect 98000 300160 98052 300212
rect 63316 300092 63368 300144
rect 132684 300092 132736 300144
rect 102324 299752 102376 299804
rect 213276 299752 213328 299804
rect 89812 299684 89864 299736
rect 232596 299684 232648 299736
rect 80612 299616 80664 299668
rect 238024 299616 238076 299668
rect 97356 299548 97408 299600
rect 333244 299548 333296 299600
rect 88432 299480 88484 299532
rect 335360 299480 335412 299532
rect 83464 298800 83516 298852
rect 127164 298800 127216 298852
rect 60464 298732 60516 298784
rect 105544 298732 105596 298784
rect 84200 298392 84252 298444
rect 144184 298392 144236 298444
rect 87420 298324 87472 298376
rect 210516 298324 210568 298376
rect 111248 298256 111300 298308
rect 318064 298256 318116 298308
rect 111892 298188 111944 298240
rect 343732 298188 343784 298240
rect 86776 298120 86828 298172
rect 320824 298120 320876 298172
rect 117412 298052 117464 298104
rect 121552 298052 121604 298104
rect 94504 297440 94556 297492
rect 107752 297440 107804 297492
rect 98644 297372 98696 297424
rect 125876 297372 125928 297424
rect 112536 296896 112588 296948
rect 202236 296896 202288 296948
rect 67548 296828 67600 296880
rect 207664 296828 207716 296880
rect 3424 296760 3476 296812
rect 100024 296760 100076 296812
rect 108672 296760 108724 296812
rect 114652 296760 114704 296812
rect 117044 296760 117096 296812
rect 342352 296760 342404 296812
rect 99012 296692 99064 296744
rect 358820 296692 358872 296744
rect 11704 295944 11756 295996
rect 71320 295944 71372 295996
rect 72424 295944 72476 295996
rect 82912 295672 82964 295724
rect 141424 295672 141476 295724
rect 40684 295604 40736 295656
rect 117320 295604 117372 295656
rect 118332 295604 118384 295656
rect 93216 295536 93268 295588
rect 203524 295536 203576 295588
rect 83556 295468 83608 295520
rect 247684 295468 247736 295520
rect 65984 295400 66036 295452
rect 240784 295400 240836 295452
rect 109316 295332 109368 295384
rect 319536 295332 319588 295384
rect 101404 295264 101456 295316
rect 104808 295264 104860 295316
rect 92756 295128 92808 295180
rect 94412 295128 94464 295180
rect 85488 294924 85540 294976
rect 87604 294924 87656 294976
rect 66168 294720 66220 294772
rect 78404 294720 78456 294772
rect 14464 294584 14516 294636
rect 53656 294584 53708 294636
rect 79048 294652 79100 294704
rect 62028 294584 62080 294636
rect 91284 294584 91336 294636
rect 70032 294380 70084 294432
rect 117964 294380 118016 294432
rect 73160 294312 73212 294364
rect 73620 294312 73672 294364
rect 88340 294312 88392 294364
rect 89076 294312 89128 294364
rect 93952 294312 94004 294364
rect 94780 294312 94832 294364
rect 100024 294312 100076 294364
rect 101588 294312 101640 294364
rect 106280 294312 106332 294364
rect 107108 294312 107160 294364
rect 110328 294312 110380 294364
rect 119804 294312 119856 294364
rect 88064 294244 88116 294296
rect 57888 294108 57940 294160
rect 96436 294176 96488 294228
rect 105452 294244 105504 294296
rect 106096 294244 106148 294296
rect 125048 294244 125100 294296
rect 114468 294176 114520 294228
rect 118976 294176 119028 294228
rect 218704 294176 218756 294228
rect 95792 294108 95844 294160
rect 195336 294108 195388 294160
rect 91928 294040 91980 294092
rect 262220 294040 262272 294092
rect 80152 293972 80204 294024
rect 92756 293972 92808 294024
rect 114376 293972 114428 294024
rect 357440 293972 357492 294024
rect 53104 293292 53156 293344
rect 56416 293292 56468 293344
rect 97080 293292 97132 293344
rect 3608 293224 3660 293276
rect 80152 293224 80204 293276
rect 114468 293224 114520 293276
rect 142804 293224 142856 293276
rect 110604 292816 110656 292868
rect 209228 292816 209280 292868
rect 117688 292748 117740 292800
rect 216128 292748 216180 292800
rect 93860 292680 93912 292732
rect 231124 292680 231176 292732
rect 99656 292612 99708 292664
rect 276112 292612 276164 292664
rect 3516 292544 3568 292596
rect 11704 292544 11756 292596
rect 68652 292544 68704 292596
rect 351920 292544 351972 292596
rect 121460 292476 121512 292528
rect 125600 292476 125652 292528
rect 103520 292068 103572 292120
rect 108304 291864 108356 291916
rect 117964 291864 118016 291916
rect 249064 291796 249116 291848
rect 249156 291252 249208 291304
rect 350632 291184 350684 291236
rect 269764 291116 269816 291168
rect 276020 291116 276072 291168
rect 121460 289892 121512 289944
rect 222936 289892 222988 289944
rect 21364 289824 21416 289876
rect 68008 289824 68060 289876
rect 121736 289824 121788 289876
rect 251824 289824 251876 289876
rect 121460 289756 121512 289808
rect 124312 289756 124364 289808
rect 119804 289076 119856 289128
rect 580264 289076 580316 289128
rect 121460 288328 121512 288380
rect 133972 288328 134024 288380
rect 135168 288328 135220 288380
rect 135168 287648 135220 287700
rect 582932 287648 582984 287700
rect 121736 287036 121788 287088
rect 345020 287036 345072 287088
rect 65984 286968 66036 287020
rect 67732 286968 67784 287020
rect 121460 286968 121512 287020
rect 127072 286968 127124 287020
rect 120908 286356 120960 286408
rect 136824 286356 136876 286408
rect 122288 286288 122340 286340
rect 328736 286288 328788 286340
rect 120816 285676 120868 285728
rect 177304 285676 177356 285728
rect 66076 285608 66128 285660
rect 68192 285608 68244 285660
rect 121736 285608 121788 285660
rect 125784 285608 125836 285660
rect 121552 284316 121604 284368
rect 311164 284316 311216 284368
rect 60648 284248 60700 284300
rect 67640 284248 67692 284300
rect 121460 284248 121512 284300
rect 128544 284248 128596 284300
rect 121460 282888 121512 282940
rect 325700 282888 325752 282940
rect 57796 282820 57848 282872
rect 67640 282820 67692 282872
rect 121460 281528 121512 281580
rect 240876 281528 240928 281580
rect 121460 280236 121512 280288
rect 227076 280236 227128 280288
rect 52184 280168 52236 280220
rect 67640 280168 67692 280220
rect 121552 280168 121604 280220
rect 247776 280168 247828 280220
rect 46756 280100 46808 280152
rect 67732 280100 67784 280152
rect 59268 280032 59320 280084
rect 67640 280032 67692 280084
rect 25504 279420 25556 279472
rect 46756 279420 46808 279472
rect 121736 279420 121788 279472
rect 255320 279420 255372 279472
rect 121460 278808 121512 278860
rect 148324 278808 148376 278860
rect 121552 278740 121604 278792
rect 312544 278740 312596 278792
rect 48044 277448 48096 277500
rect 67640 277448 67692 277500
rect 121460 277448 121512 277500
rect 315304 277448 315356 277500
rect 46848 277380 46900 277432
rect 67732 277380 67784 277432
rect 121552 277380 121604 277432
rect 322204 277380 322256 277432
rect 121460 277312 121512 277364
rect 129924 277312 129976 277364
rect 129924 276632 129976 276684
rect 144092 276632 144144 276684
rect 50804 276088 50856 276140
rect 67640 276088 67692 276140
rect 121460 276020 121512 276072
rect 338212 276020 338264 276072
rect 64604 274728 64656 274780
rect 67640 274728 67692 274780
rect 57796 274660 57848 274712
rect 67824 274660 67876 274712
rect 44088 274592 44140 274644
rect 67732 274592 67784 274644
rect 121460 274592 121512 274644
rect 124864 274592 124916 274644
rect 121644 273912 121696 273964
rect 468484 273912 468536 273964
rect 121460 273232 121512 273284
rect 214564 273232 214616 273284
rect 121552 273164 121604 273216
rect 125876 273164 125928 273216
rect 139400 273164 139452 273216
rect 580172 273164 580224 273216
rect 124956 272484 125008 272536
rect 139400 272484 139452 272536
rect 60280 271940 60332 271992
rect 67640 271940 67692 271992
rect 59268 271872 59320 271924
rect 67824 271872 67876 271924
rect 60556 271804 60608 271856
rect 67732 271804 67784 271856
rect 61752 270512 61804 270564
rect 67640 270512 67692 270564
rect 121460 270512 121512 270564
rect 252652 270512 252704 270564
rect 144092 269764 144144 269816
rect 580540 269764 580592 269816
rect 54760 269152 54812 269204
rect 67732 269152 67784 269204
rect 53656 269084 53708 269136
rect 67640 269084 67692 269136
rect 121460 269084 121512 269136
rect 233884 269084 233936 269136
rect 121552 269016 121604 269068
rect 132592 269016 132644 269068
rect 43996 268336 44048 268388
rect 67640 268336 67692 268388
rect 121644 268336 121696 268388
rect 252560 268336 252612 268388
rect 66168 268200 66220 268252
rect 68192 268200 68244 268252
rect 43444 268064 43496 268116
rect 43996 268064 44048 268116
rect 121460 267724 121512 267776
rect 339500 267724 339552 267776
rect 41328 267656 41380 267708
rect 67732 267656 67784 267708
rect 54944 267588 54996 267640
rect 67640 267588 67692 267640
rect 3332 267112 3384 267164
rect 7564 267112 7616 267164
rect 121460 266432 121512 266484
rect 334072 266432 334124 266484
rect 121552 266364 121604 266416
rect 347964 266364 348016 266416
rect 53564 266296 53616 266348
rect 67640 266296 67692 266348
rect 125048 265616 125100 265668
rect 580448 265616 580500 265668
rect 121460 265004 121512 265056
rect 308496 265004 308548 265056
rect 56232 264936 56284 264988
rect 67732 264936 67784 264988
rect 121552 264936 121604 264988
rect 346492 264936 346544 264988
rect 48136 264868 48188 264920
rect 67640 264868 67692 264920
rect 121460 264868 121512 264920
rect 125692 264868 125744 264920
rect 18604 264188 18656 264240
rect 48136 264188 48188 264240
rect 49516 263576 49568 263628
rect 67732 263576 67784 263628
rect 121552 263576 121604 263628
rect 233976 263576 234028 263628
rect 50896 263508 50948 263560
rect 67640 263508 67692 263560
rect 121460 263508 121512 263560
rect 123116 263508 123168 263560
rect 59084 262216 59136 262268
rect 67640 262216 67692 262268
rect 121460 262216 121512 262268
rect 338396 262216 338448 262268
rect 54852 260924 54904 260976
rect 67640 260924 67692 260976
rect 53564 260856 53616 260908
rect 67732 260856 67784 260908
rect 121552 260856 121604 260908
rect 307116 260856 307168 260908
rect 61936 260788 61988 260840
rect 67640 260788 67692 260840
rect 121460 260788 121512 260840
rect 142160 260788 142212 260840
rect 143448 260788 143500 260840
rect 143448 260108 143500 260160
rect 464344 260108 464396 260160
rect 61384 259428 61436 259480
rect 67640 259428 67692 259480
rect 121460 259428 121512 259480
rect 235264 259428 235316 259480
rect 121552 259360 121604 259412
rect 132500 259360 132552 259412
rect 273904 259360 273956 259412
rect 579896 259360 579948 259412
rect 60372 258136 60424 258188
rect 67640 258136 67692 258188
rect 56416 258068 56468 258120
rect 67732 258068 67784 258120
rect 121644 258068 121696 258120
rect 347872 258068 347924 258120
rect 34336 258000 34388 258052
rect 67640 258000 67692 258052
rect 121460 258000 121512 258052
rect 129004 258000 129056 258052
rect 63316 257388 63368 257440
rect 68376 257388 68428 257440
rect 4804 257320 4856 257372
rect 34336 257320 34388 257372
rect 60648 257320 60700 257372
rect 68284 257320 68336 257372
rect 63224 256708 63276 256760
rect 67640 256708 67692 256760
rect 121552 256708 121604 256760
rect 220084 256708 220136 256760
rect 121460 256640 121512 256692
rect 129832 256640 129884 256692
rect 121552 256572 121604 256624
rect 126980 256572 127032 256624
rect 120908 255960 120960 256012
rect 580356 255960 580408 256012
rect 3148 255212 3200 255264
rect 34888 255212 34940 255264
rect 55128 255212 55180 255264
rect 67640 255212 67692 255264
rect 56324 254600 56376 254652
rect 61660 254600 61712 254652
rect 67640 254600 67692 254652
rect 34888 254532 34940 254584
rect 35808 254532 35860 254584
rect 58624 254532 58676 254584
rect 121460 253988 121512 254040
rect 246396 253988 246448 254040
rect 121552 253920 121604 253972
rect 314016 253920 314068 253972
rect 54484 253852 54536 253904
rect 56508 253852 56560 253904
rect 67640 253852 67692 253904
rect 121552 252628 121604 252680
rect 263600 252628 263652 252680
rect 64512 252560 64564 252612
rect 67640 252560 67692 252612
rect 121460 252560 121512 252612
rect 350724 252560 350776 252612
rect 64696 251268 64748 251320
rect 67732 251268 67784 251320
rect 56508 251200 56560 251252
rect 67640 251200 67692 251252
rect 121460 251200 121512 251252
rect 331312 251200 331364 251252
rect 120448 250996 120500 251048
rect 123024 250996 123076 251048
rect 65892 249840 65944 249892
rect 67640 249840 67692 249892
rect 57612 249772 57664 249824
rect 67732 249772 67784 249824
rect 121552 249772 121604 249824
rect 238116 249772 238168 249824
rect 49608 249704 49660 249756
rect 67640 249704 67692 249756
rect 121460 249704 121512 249756
rect 140872 249704 140924 249756
rect 59176 249636 59228 249688
rect 61384 249636 61436 249688
rect 120724 249500 120776 249552
rect 121460 249500 121512 249552
rect 66076 248616 66128 248668
rect 68100 248616 68152 248668
rect 121552 248412 121604 248464
rect 210424 248412 210476 248464
rect 121460 248344 121512 248396
rect 121644 248344 121696 248396
rect 147680 248344 147732 248396
rect 121736 248276 121788 248328
rect 177304 247664 177356 247716
rect 580356 247664 580408 247716
rect 62028 247120 62080 247172
rect 67732 247120 67784 247172
rect 61936 247052 61988 247104
rect 67640 247052 67692 247104
rect 121460 247052 121512 247104
rect 266360 247052 266412 247104
rect 121552 245692 121604 245744
rect 224316 245692 224368 245744
rect 121460 245624 121512 245676
rect 231216 245624 231268 245676
rect 61844 245556 61896 245608
rect 67640 245556 67692 245608
rect 65984 244264 66036 244316
rect 68100 244264 68152 244316
rect 342444 244264 342496 244316
rect 580172 244264 580224 244316
rect 11704 244196 11756 244248
rect 39856 244196 39908 244248
rect 67640 244196 67692 244248
rect 121460 244196 121512 244248
rect 134064 244196 134116 244248
rect 121644 243516 121696 243568
rect 321560 243516 321612 243568
rect 121552 242904 121604 242956
rect 335544 242904 335596 242956
rect 121460 242836 121512 242888
rect 132684 242836 132736 242888
rect 342444 242836 342496 242888
rect 121552 242768 121604 242820
rect 128452 242768 128504 242820
rect 63408 241476 63460 241528
rect 67640 241476 67692 241528
rect 121460 241476 121512 241528
rect 249800 241476 249852 241528
rect 121552 240728 121604 240780
rect 135260 240728 135312 240780
rect 3056 240116 3108 240168
rect 11152 240116 11204 240168
rect 119896 240116 119948 240168
rect 329840 240116 329892 240168
rect 65892 239912 65944 239964
rect 72516 239912 72568 239964
rect 75920 239776 75972 239828
rect 77104 239776 77156 239828
rect 78680 239776 78732 239828
rect 79680 239776 79732 239828
rect 86960 239776 87012 239828
rect 88052 239776 88104 239828
rect 89720 239776 89772 239828
rect 90628 239776 90680 239828
rect 100760 239776 100812 239828
rect 101576 239776 101628 239828
rect 103612 239776 103664 239828
rect 104796 239776 104848 239828
rect 104900 239776 104952 239828
rect 106084 239776 106136 239828
rect 107660 239776 107712 239828
rect 108660 239776 108712 239828
rect 114560 239776 114612 239828
rect 115744 239776 115796 239828
rect 121460 239708 121512 239760
rect 124864 239708 124916 239760
rect 69756 239504 69808 239556
rect 83556 239504 83608 239556
rect 64512 239436 64564 239488
rect 339592 239436 339644 239488
rect 63224 239368 63276 239420
rect 342444 239368 342496 239420
rect 84292 239300 84344 239352
rect 85488 239300 85540 239352
rect 99012 238960 99064 239012
rect 131120 238960 131172 239012
rect 115112 238892 115164 238944
rect 124220 238892 124272 238944
rect 114468 238824 114520 238876
rect 127164 238824 127216 238876
rect 52368 238756 52420 238808
rect 95792 238756 95844 238808
rect 7564 238688 7616 238740
rect 57704 238688 57756 238740
rect 86776 238688 86828 238740
rect 89352 238688 89404 238740
rect 129740 238688 129792 238740
rect 48228 238620 48280 238672
rect 82268 238620 82320 238672
rect 91928 238620 91980 238672
rect 120908 238620 120960 238672
rect 63132 238552 63184 238604
rect 72608 238552 72660 238604
rect 118332 238552 118384 238604
rect 136732 238552 136784 238604
rect 106740 238484 106792 238536
rect 121460 238484 121512 238536
rect 102876 238144 102928 238196
rect 106924 238144 106976 238196
rect 82912 238076 82964 238128
rect 88984 238076 89036 238128
rect 96436 238076 96488 238128
rect 184204 238076 184256 238128
rect 68836 238008 68888 238060
rect 327172 238008 327224 238060
rect 71320 237464 71372 237516
rect 75184 237464 75236 237516
rect 69940 237396 69992 237448
rect 72424 237396 72476 237448
rect 75828 237328 75880 237380
rect 143540 237328 143592 237380
rect 68928 236648 68980 236700
rect 286324 236648 286376 236700
rect 324964 236648 325016 236700
rect 347780 236648 347832 236700
rect 11152 235900 11204 235952
rect 37096 235900 37148 235952
rect 103520 235900 103572 235952
rect 117688 235900 117740 235952
rect 133880 235900 133932 235952
rect 135168 235900 135220 235952
rect 58624 235832 58676 235884
rect 112536 235832 112588 235884
rect 53748 235764 53800 235816
rect 107384 235764 107436 235816
rect 52276 235696 52328 235748
rect 76564 235696 76616 235748
rect 81624 235696 81676 235748
rect 120816 235696 120868 235748
rect 91284 235628 91336 235680
rect 124956 235628 125008 235680
rect 135168 235220 135220 235272
rect 180156 235220 180208 235272
rect 45468 234540 45520 234592
rect 109040 234540 109092 234592
rect 110604 234540 110656 234592
rect 111064 234540 111116 234592
rect 136640 234540 136692 234592
rect 88984 234472 89036 234524
rect 128360 234472 128412 234524
rect 109040 234132 109092 234184
rect 109960 234132 110012 234184
rect 80336 233928 80388 233980
rect 320916 233928 320968 233980
rect 128360 233860 128412 233912
rect 582748 233860 582800 233912
rect 84108 231820 84160 231872
rect 84844 231820 84896 231872
rect 64604 231140 64656 231192
rect 133144 231140 133196 231192
rect 78312 231072 78364 231124
rect 267740 231072 267792 231124
rect 60188 230392 60240 230444
rect 60464 230392 60516 230444
rect 83372 230392 83424 230444
rect 17224 229712 17276 229764
rect 60188 229712 60240 229764
rect 72516 229712 72568 229764
rect 336740 229712 336792 229764
rect 97632 228420 97684 228472
rect 333980 228420 334032 228472
rect 88340 228352 88392 228404
rect 353392 228352 353444 228404
rect 63408 226992 63460 227044
rect 214656 226992 214708 227044
rect 3608 225564 3660 225616
rect 120080 225564 120132 225616
rect 78772 224272 78824 224324
rect 228364 224272 228416 224324
rect 95056 224204 95108 224256
rect 345112 224204 345164 224256
rect 75184 221484 75236 221536
rect 242164 221484 242216 221536
rect 56232 221416 56284 221468
rect 340880 221416 340932 221468
rect 114560 220124 114612 220176
rect 311256 220124 311308 220176
rect 46848 220056 46900 220108
rect 296076 220056 296128 220108
rect 110420 218764 110472 218816
rect 256976 218764 257028 218816
rect 103612 218696 103664 218748
rect 325792 218696 325844 218748
rect 82084 217268 82136 217320
rect 300216 217268 300268 217320
rect 99472 215976 99524 216028
rect 253940 215976 253992 216028
rect 93952 215908 94004 215960
rect 322940 215908 322992 215960
rect 3332 215228 3384 215280
rect 18604 215228 18656 215280
rect 56416 214616 56468 214668
rect 280160 214616 280212 214668
rect 103704 214548 103756 214600
rect 352104 214548 352156 214600
rect 89812 213324 89864 213376
rect 254124 213324 254176 213376
rect 87052 213256 87104 213308
rect 327080 213256 327132 213308
rect 54852 213188 54904 213240
rect 316684 213188 316736 213240
rect 104992 211760 105044 211812
rect 331496 211760 331548 211812
rect 61936 210468 61988 210520
rect 236644 210468 236696 210520
rect 83464 210400 83516 210452
rect 335452 210400 335504 210452
rect 100852 209176 100904 209228
rect 254032 209176 254084 209228
rect 48044 209108 48096 209160
rect 270500 209108 270552 209160
rect 113180 209040 113232 209092
rect 338304 209040 338356 209092
rect 86960 207680 87012 207732
rect 252836 207680 252888 207732
rect 74632 207612 74684 207664
rect 278872 207612 278924 207664
rect 111800 206252 111852 206304
rect 255412 206252 255464 206304
rect 89720 204960 89772 205012
rect 281632 204960 281684 205012
rect 59084 204892 59136 204944
rect 259460 204892 259512 204944
rect 50804 203532 50856 203584
rect 263784 203532 263836 203584
rect 106924 202240 106976 202292
rect 239404 202240 239456 202292
rect 100760 202172 100812 202224
rect 252744 202172 252796 202224
rect 72424 202104 72476 202156
rect 343916 202104 343968 202156
rect 93860 200880 93912 200932
rect 255504 200880 255556 200932
rect 96620 200812 96672 200864
rect 260840 200812 260892 200864
rect 107752 200744 107804 200796
rect 328644 200744 328696 200796
rect 133144 199520 133196 199572
rect 265072 199520 265124 199572
rect 115940 199452 115992 199504
rect 270684 199452 270736 199504
rect 77300 199384 77352 199436
rect 329932 199384 329984 199436
rect 251824 198160 251876 198212
rect 274824 198160 274876 198212
rect 60280 198092 60332 198144
rect 272064 198092 272116 198144
rect 92572 198024 92624 198076
rect 330024 198024 330076 198076
rect 76564 197956 76616 198008
rect 582840 197956 582892 198008
rect 92480 196732 92532 196784
rect 261024 196732 261076 196784
rect 69020 196664 69072 196716
rect 251180 196664 251232 196716
rect 107660 196596 107712 196648
rect 328552 196596 328604 196648
rect 54760 195372 54812 195424
rect 269212 195372 269264 195424
rect 124864 195304 124916 195356
rect 345204 195304 345256 195356
rect 86224 195236 86276 195288
rect 582656 195236 582708 195288
rect 247776 194012 247828 194064
rect 340972 194012 341024 194064
rect 142804 193944 142856 193996
rect 259736 193944 259788 193996
rect 57612 193876 57664 193928
rect 273352 193876 273404 193928
rect 78680 193808 78732 193860
rect 335636 193808 335688 193860
rect 152464 192720 152516 192772
rect 200764 192720 200816 192772
rect 146944 192652 146996 192704
rect 209136 192652 209188 192704
rect 199384 192584 199436 192636
rect 280252 192584 280304 192636
rect 84292 192516 84344 192568
rect 254216 192516 254268 192568
rect 70400 192448 70452 192500
rect 321744 192448 321796 192500
rect 148324 191292 148376 191344
rect 239496 191292 239548 191344
rect 246304 191292 246356 191344
rect 277492 191292 277544 191344
rect 192484 191224 192536 191276
rect 331404 191224 331456 191276
rect 59268 191156 59320 191208
rect 256792 191156 256844 191208
rect 62028 191088 62080 191140
rect 262312 191088 262364 191140
rect 213276 189864 213328 189916
rect 281724 189864 281776 189916
rect 144184 189796 144236 189848
rect 242256 189796 242308 189848
rect 56508 189728 56560 189780
rect 199476 189728 199528 189780
rect 249156 189728 249208 189780
rect 336832 189728 336884 189780
rect 107568 189048 107620 189100
rect 188436 189048 188488 189100
rect 209228 188640 209280 188692
rect 261116 188640 261168 188692
rect 202236 188572 202288 188624
rect 267924 188572 267976 188624
rect 15844 188504 15896 188556
rect 109040 188504 109092 188556
rect 141424 188504 141476 188556
rect 262404 188504 262456 188556
rect 69204 188436 69256 188488
rect 319628 188436 319680 188488
rect 69112 188368 69164 188420
rect 341156 188368 341208 188420
rect 57796 188300 57848 188352
rect 334256 188300 334308 188352
rect 129648 187756 129700 187808
rect 177304 187756 177356 187808
rect 104808 187688 104860 187740
rect 173256 187688 173308 187740
rect 203524 187008 203576 187060
rect 276204 187008 276256 187060
rect 73252 186940 73304 186992
rect 323124 186940 323176 186992
rect 100668 186464 100720 186516
rect 169116 186464 169168 186516
rect 99288 186396 99340 186448
rect 171784 186396 171836 186448
rect 119988 186328 120040 186380
rect 214748 186328 214800 186380
rect 151084 185920 151136 185972
rect 187056 185920 187108 185972
rect 232596 185920 232648 185972
rect 266452 185920 266504 185972
rect 65984 185852 66036 185904
rect 274732 185852 274784 185904
rect 99380 185784 99432 185836
rect 325976 185784 326028 185836
rect 104900 185716 104952 185768
rect 339684 185716 339736 185768
rect 80060 185648 80112 185700
rect 327356 185648 327408 185700
rect 67456 185580 67508 185632
rect 324320 185580 324372 185632
rect 214656 184356 214708 184408
rect 270592 184356 270644 184408
rect 67548 184288 67600 184340
rect 251272 184288 251324 184340
rect 73160 184220 73212 184272
rect 323216 184220 323268 184272
rect 64696 184152 64748 184204
rect 341064 184152 341116 184204
rect 128268 183608 128320 183660
rect 166540 183608 166592 183660
rect 114468 183540 114520 183592
rect 169300 183540 169352 183592
rect 224224 183132 224276 183184
rect 258264 183132 258316 183184
rect 226984 183064 227036 183116
rect 263876 183064 263928 183116
rect 155224 182996 155276 183048
rect 193864 182996 193916 183048
rect 222844 182996 222896 183048
rect 266544 182996 266596 183048
rect 311164 182996 311216 183048
rect 332784 182996 332836 183048
rect 63316 182928 63368 182980
rect 271972 182928 272024 182980
rect 307116 182928 307168 182980
rect 334164 182928 334216 182980
rect 84200 182860 84252 182912
rect 325884 182860 325936 182912
rect 75920 182792 75972 182844
rect 321652 182792 321704 182844
rect 116952 182248 117004 182300
rect 170588 182248 170640 182300
rect 110696 182180 110748 182232
rect 167644 182180 167696 182232
rect 231216 181704 231268 181756
rect 258080 181704 258132 181756
rect 238024 181636 238076 181688
rect 264980 181636 265032 181688
rect 122104 181568 122156 181620
rect 171140 181568 171192 181620
rect 207664 181568 207716 181620
rect 273536 181568 273588 181620
rect 59176 181500 59228 181552
rect 336924 181500 336976 181552
rect 53564 181432 53616 181484
rect 345296 181432 345348 181484
rect 120908 180956 120960 181008
rect 167736 180956 167788 181008
rect 115848 180888 115900 180940
rect 166448 180888 166500 180940
rect 130752 180820 130804 180872
rect 214656 180820 214708 180872
rect 239404 180412 239456 180464
rect 258356 180412 258408 180464
rect 233976 180344 234028 180396
rect 265256 180344 265308 180396
rect 166264 180276 166316 180328
rect 182824 180276 182876 180328
rect 222936 180276 222988 180328
rect 263692 180276 263744 180328
rect 160744 180208 160796 180260
rect 192484 180208 192536 180260
rect 220084 180208 220136 180260
rect 267832 180208 267884 180260
rect 66076 180140 66128 180192
rect 273444 180140 273496 180192
rect 300124 180140 300176 180192
rect 332600 180140 332652 180192
rect 71872 180072 71924 180124
rect 327264 180072 327316 180124
rect 125416 179460 125468 179512
rect 167920 179460 167972 179512
rect 112168 179392 112220 179444
rect 170496 179392 170548 179444
rect 235264 178916 235316 178968
rect 265164 178916 265216 178968
rect 227076 178848 227128 178900
rect 259552 178848 259604 178900
rect 214564 178780 214616 178832
rect 249340 178780 249392 178832
rect 315304 178780 315356 178832
rect 339776 178780 339828 178832
rect 66168 178712 66220 178764
rect 251364 178712 251416 178764
rect 311256 178712 311308 178764
rect 342536 178712 342588 178764
rect 102140 178644 102192 178696
rect 346584 178644 346636 178696
rect 133144 178236 133196 178288
rect 164884 178236 164936 178288
rect 148232 178168 148284 178220
rect 181444 178168 181496 178220
rect 123300 178100 123352 178152
rect 166356 178100 166408 178152
rect 110052 178032 110104 178084
rect 170404 178032 170456 178084
rect 272616 178032 272668 178084
rect 316040 178032 316092 178084
rect 242164 177964 242216 178016
rect 249892 177964 249944 178016
rect 247684 177556 247736 177608
rect 258172 177556 258224 177608
rect 319536 177556 319588 177608
rect 330116 177556 330168 177608
rect 233884 177488 233936 177540
rect 260932 177488 260984 177540
rect 319628 177488 319680 177540
rect 331220 177488 331272 177540
rect 228364 177420 228416 177472
rect 259644 177420 259696 177472
rect 314016 177420 314068 177472
rect 332692 177420 332744 177472
rect 224316 177352 224368 177404
rect 262496 177352 262548 177404
rect 307024 177352 307076 177404
rect 350540 177352 350592 177404
rect 184204 177284 184256 177336
rect 324412 177284 324464 177336
rect 333244 177284 333296 177336
rect 338120 177284 338172 177336
rect 134432 177012 134484 177064
rect 165436 177012 165488 177064
rect 103336 176944 103388 176996
rect 169208 176944 169260 176996
rect 108120 176876 108172 176928
rect 184848 176876 184900 176928
rect 136088 176808 136140 176860
rect 213920 176808 213972 176860
rect 125876 176740 125928 176792
rect 214932 176740 214984 176792
rect 102048 176672 102100 176724
rect 202236 176672 202288 176724
rect 132040 176264 132092 176316
rect 165528 176264 165580 176316
rect 158904 176196 158956 176248
rect 198096 176196 198148 176248
rect 238116 176196 238168 176248
rect 249248 176196 249300 176248
rect 118424 176128 118476 176180
rect 166264 176128 166316 176180
rect 239496 176128 239548 176180
rect 249064 176128 249116 176180
rect 319444 176128 319496 176180
rect 326160 176128 326212 176180
rect 121920 176060 121972 176112
rect 170680 176060 170732 176112
rect 246396 176060 246448 176112
rect 255596 176060 255648 176112
rect 312544 176060 312596 176112
rect 321468 176060 321520 176112
rect 100760 175992 100812 176044
rect 184204 175992 184256 176044
rect 184848 175992 184900 176044
rect 214564 175992 214616 176044
rect 316684 175992 316736 176044
rect 332876 175992 332928 176044
rect 11704 175924 11756 175976
rect 111064 175924 111116 175976
rect 127072 175924 127124 175976
rect 211896 175924 211948 175976
rect 236644 175924 236696 175976
rect 256884 175924 256936 175976
rect 318064 175924 318116 175976
rect 337016 175924 337068 175976
rect 165436 175176 165488 175228
rect 213920 175176 213972 175228
rect 164884 175108 164936 175160
rect 214012 175108 214064 175160
rect 291936 174020 291988 174072
rect 307668 174020 307720 174072
rect 289176 173952 289228 174004
rect 307484 173952 307536 174004
rect 269764 173884 269816 173936
rect 307576 173884 307628 173936
rect 165528 173816 165580 173868
rect 213920 173816 213972 173868
rect 252468 173816 252520 173868
rect 263784 173816 263836 173868
rect 324320 173816 324372 173868
rect 326160 173816 326212 173868
rect 295984 172660 296036 172712
rect 307484 172660 307536 172712
rect 289084 172592 289136 172644
rect 307576 172592 307628 172644
rect 267004 172524 267056 172576
rect 307668 172524 307720 172576
rect 166540 172456 166592 172508
rect 214012 172456 214064 172508
rect 177304 172388 177356 172440
rect 213920 172388 213972 172440
rect 252468 172320 252520 172372
rect 266360 172320 266412 172372
rect 296076 171232 296128 171284
rect 306564 171232 306616 171284
rect 268384 171164 268436 171216
rect 307576 171164 307628 171216
rect 264428 171096 264480 171148
rect 307668 171096 307720 171148
rect 211896 171028 211948 171080
rect 214472 171028 214524 171080
rect 252376 171028 252428 171080
rect 265072 171028 265124 171080
rect 324320 171028 324372 171080
rect 338120 171028 338172 171080
rect 252284 170824 252336 170876
rect 256884 170824 256936 170876
rect 252468 170756 252520 170808
rect 258264 170756 258316 170808
rect 300124 169872 300176 169924
rect 307668 169872 307720 169924
rect 286416 169804 286468 169856
rect 307300 169804 307352 169856
rect 259092 169736 259144 169788
rect 262220 169736 262272 169788
rect 275376 169736 275428 169788
rect 307484 169736 307536 169788
rect 166356 169668 166408 169720
rect 214012 169668 214064 169720
rect 252376 169668 252428 169720
rect 260840 169668 260892 169720
rect 324320 169668 324372 169720
rect 345296 169668 345348 169720
rect 167920 169600 167972 169652
rect 213920 169600 213972 169652
rect 252468 169056 252520 169108
rect 258356 169056 258408 169108
rect 252468 168648 252520 168700
rect 259736 168648 259788 168700
rect 290464 168512 290516 168564
rect 307116 168512 307168 168564
rect 271328 168444 271380 168496
rect 307668 168444 307720 168496
rect 262864 168376 262916 168428
rect 307576 168376 307628 168428
rect 167736 168308 167788 168360
rect 214012 168308 214064 168360
rect 252376 168308 252428 168360
rect 263600 168308 263652 168360
rect 324320 168308 324372 168360
rect 339592 168308 339644 168360
rect 170680 168240 170732 168292
rect 213920 168240 213972 168292
rect 252468 168240 252520 168292
rect 262404 168240 262456 168292
rect 324412 168240 324464 168292
rect 331220 168240 331272 168292
rect 252468 167220 252520 167272
rect 259092 167220 259144 167272
rect 283748 167152 283800 167204
rect 307484 167152 307536 167204
rect 281080 167084 281132 167136
rect 307668 167084 307720 167136
rect 276664 167016 276716 167068
rect 307300 167016 307352 167068
rect 166264 166948 166316 167000
rect 214012 166948 214064 167000
rect 252376 166948 252428 167000
rect 261024 166948 261076 167000
rect 324320 166948 324372 167000
rect 346676 166948 346728 167000
rect 464344 166948 464396 167000
rect 580172 166948 580224 167000
rect 170588 166880 170640 166932
rect 213920 166880 213972 166932
rect 252468 166812 252520 166864
rect 259460 166812 259512 166864
rect 302884 165724 302936 165776
rect 307116 165724 307168 165776
rect 278228 165656 278280 165708
rect 307576 165656 307628 165708
rect 260196 165588 260248 165640
rect 307668 165588 307720 165640
rect 166448 165520 166500 165572
rect 213920 165520 213972 165572
rect 252376 165520 252428 165572
rect 270500 165520 270552 165572
rect 324412 165520 324464 165572
rect 346584 165520 346636 165572
rect 169300 165452 169352 165504
rect 214012 165452 214064 165504
rect 252468 165452 252520 165504
rect 261116 165452 261168 165504
rect 324320 165452 324372 165504
rect 343916 165452 343968 165504
rect 251364 165384 251416 165436
rect 254124 165384 254176 165436
rect 269856 164840 269908 164892
rect 307392 164840 307444 164892
rect 305736 164296 305788 164348
rect 307116 164296 307168 164348
rect 287980 164228 288032 164280
rect 307668 164228 307720 164280
rect 3240 164160 3292 164212
rect 14464 164160 14516 164212
rect 170496 164160 170548 164212
rect 213920 164160 213972 164212
rect 252376 164160 252428 164212
rect 266544 164160 266596 164212
rect 324412 164160 324464 164212
rect 336924 164160 336976 164212
rect 252284 164092 252336 164144
rect 265256 164092 265308 164144
rect 324320 164092 324372 164144
rect 332876 164092 332928 164144
rect 252468 164024 252520 164076
rect 263876 164024 263928 164076
rect 301504 163004 301556 163056
rect 307576 163004 307628 163056
rect 271236 162936 271288 162988
rect 306748 162936 306800 162988
rect 257528 162868 257580 162920
rect 307668 162868 307720 162920
rect 167644 162800 167696 162852
rect 213920 162800 213972 162852
rect 324412 162800 324464 162852
rect 335544 162800 335596 162852
rect 170404 162732 170456 162784
rect 214012 162732 214064 162784
rect 252468 162732 252520 162784
rect 267740 162732 267792 162784
rect 324320 162732 324372 162784
rect 330116 162732 330168 162784
rect 297456 161576 297508 161628
rect 307484 161576 307536 161628
rect 264244 161508 264296 161560
rect 307576 161508 307628 161560
rect 258908 161440 258960 161492
rect 307668 161440 307720 161492
rect 188436 161372 188488 161424
rect 213920 161372 213972 161424
rect 252376 161372 252428 161424
rect 270684 161372 270736 161424
rect 324320 161372 324372 161424
rect 337016 161372 337068 161424
rect 324412 161304 324464 161356
rect 332784 161304 332836 161356
rect 252008 160964 252060 161016
rect 255320 160964 255372 161016
rect 252468 160760 252520 160812
rect 258172 160760 258224 160812
rect 167828 160692 167880 160744
rect 214656 160692 214708 160744
rect 291844 160216 291896 160268
rect 307668 160216 307720 160268
rect 265624 160148 265676 160200
rect 306564 160148 306616 160200
rect 258724 160080 258776 160132
rect 307576 160080 307628 160132
rect 173256 160012 173308 160064
rect 213920 160012 213972 160064
rect 252468 160012 252520 160064
rect 274824 160012 274876 160064
rect 298836 159332 298888 159384
rect 307208 159332 307260 159384
rect 262956 158788 263008 158840
rect 307576 158788 307628 158840
rect 254584 158720 254636 158772
rect 307668 158720 307720 158772
rect 169208 158652 169260 158704
rect 213920 158652 213972 158704
rect 252468 158652 252520 158704
rect 276204 158652 276256 158704
rect 324412 158652 324464 158704
rect 350632 158652 350684 158704
rect 202236 158584 202288 158636
rect 214012 158584 214064 158636
rect 324320 158584 324372 158636
rect 334072 158584 334124 158636
rect 293408 157496 293460 157548
rect 307668 157496 307720 157548
rect 264336 157428 264388 157480
rect 306932 157428 306984 157480
rect 258816 157360 258868 157412
rect 307576 157360 307628 157412
rect 169116 157292 169168 157344
rect 214012 157292 214064 157344
rect 252376 157292 252428 157344
rect 272064 157292 272116 157344
rect 184204 157224 184256 157276
rect 213920 157224 213972 157276
rect 252468 157224 252520 157276
rect 265164 157224 265216 157276
rect 324320 157224 324372 157276
rect 349344 157224 349396 157276
rect 324320 156816 324372 156868
rect 325976 156816 326028 156868
rect 300768 156068 300820 156120
rect 307668 156068 307720 156120
rect 268476 156000 268528 156052
rect 307484 156000 307536 156052
rect 260104 155932 260156 155984
rect 307576 155932 307628 155984
rect 171784 155864 171836 155916
rect 213920 155864 213972 155916
rect 252468 155864 252520 155916
rect 254032 155864 254084 155916
rect 324412 155864 324464 155916
rect 341156 155864 341208 155916
rect 251548 155796 251600 155848
rect 254216 155796 254268 155848
rect 324320 155796 324372 155848
rect 339776 155796 339828 155848
rect 252468 155728 252520 155780
rect 266452 155728 266504 155780
rect 282460 155184 282512 155236
rect 307392 155184 307444 155236
rect 267096 154640 267148 154692
rect 306564 154640 306616 154692
rect 254860 154572 254912 154624
rect 307668 154572 307720 154624
rect 324320 154504 324372 154556
rect 353392 154504 353444 154556
rect 252468 154436 252520 154488
rect 269212 154436 269264 154488
rect 251824 153824 251876 153876
rect 300768 153824 300820 153876
rect 324320 153416 324372 153468
rect 327356 153416 327408 153468
rect 300400 153348 300452 153400
rect 307576 153348 307628 153400
rect 178868 153280 178920 153332
rect 214012 153280 214064 153332
rect 297640 153280 297692 153332
rect 307668 153280 307720 153332
rect 175924 153212 175976 153264
rect 213920 153212 213972 153264
rect 254768 153212 254820 153264
rect 306564 153212 306616 153264
rect 252376 153144 252428 153196
rect 273536 153144 273588 153196
rect 324412 153144 324464 153196
rect 350724 153144 350776 153196
rect 252468 153076 252520 153128
rect 267924 153076 267976 153128
rect 296168 151920 296220 151972
rect 306564 151920 306616 151972
rect 184296 151852 184348 151904
rect 213920 151852 213972 151904
rect 272800 151852 272852 151904
rect 307668 151852 307720 151904
rect 177304 151784 177356 151836
rect 214012 151784 214064 151836
rect 256148 151784 256200 151836
rect 307484 151784 307536 151836
rect 252468 151716 252520 151768
rect 281632 151716 281684 151768
rect 324320 151716 324372 151768
rect 328644 151716 328696 151768
rect 252376 151648 252428 151700
rect 255412 151648 255464 151700
rect 251364 151444 251416 151496
rect 253940 151444 253992 151496
rect 300308 150560 300360 150612
rect 307668 150560 307720 150612
rect 273996 150492 274048 150544
rect 307484 150492 307536 150544
rect 199568 150424 199620 150476
rect 213920 150424 213972 150476
rect 256056 150424 256108 150476
rect 307576 150424 307628 150476
rect 3516 150356 3568 150408
rect 21364 150356 21416 150408
rect 181444 150356 181496 150408
rect 214012 150356 214064 150408
rect 252468 150356 252520 150408
rect 277492 150356 277544 150408
rect 324320 150356 324372 150408
rect 334256 150356 334308 150408
rect 252100 150288 252152 150340
rect 255504 150288 255556 150340
rect 324412 150288 324464 150340
rect 331312 150288 331364 150340
rect 252284 150220 252336 150272
rect 255596 150220 255648 150272
rect 275468 149676 275520 149728
rect 307208 149676 307260 149728
rect 255320 149336 255372 149388
rect 258080 149336 258132 149388
rect 297732 149132 297784 149184
rect 307484 149132 307536 149184
rect 254676 149064 254728 149116
rect 306564 149064 306616 149116
rect 198096 148996 198148 149048
rect 213920 148996 213972 149048
rect 252376 148996 252428 149048
rect 280252 148996 280304 149048
rect 252468 148928 252520 148980
rect 278872 148928 278924 148980
rect 324320 148928 324372 148980
rect 347964 148928 348016 148980
rect 252284 148860 252336 148912
rect 256792 148860 256844 148912
rect 259000 148316 259052 148368
rect 306656 148316 306708 148368
rect 257344 147772 257396 147824
rect 307668 147772 307720 147824
rect 167644 147636 167696 147688
rect 213920 147636 213972 147688
rect 304356 147636 304408 147688
rect 307300 147636 307352 147688
rect 324320 147568 324372 147620
rect 335360 147568 335412 147620
rect 252468 147500 252520 147552
rect 273352 147500 273404 147552
rect 252192 146888 252244 146940
rect 260932 146888 260984 146940
rect 301780 146616 301832 146668
rect 307576 146616 307628 146668
rect 210608 146344 210660 146396
rect 214012 146344 214064 146396
rect 261484 146344 261536 146396
rect 307300 146344 307352 146396
rect 174544 146276 174596 146328
rect 213920 146276 213972 146328
rect 256240 146276 256292 146328
rect 306932 146276 306984 146328
rect 252468 146208 252520 146260
rect 280160 146208 280212 146260
rect 324320 146208 324372 146260
rect 342352 146208 342404 146260
rect 252376 146140 252428 146192
rect 270592 146140 270644 146192
rect 252284 146072 252336 146124
rect 259644 146072 259696 146124
rect 324320 145664 324372 145716
rect 327172 145664 327224 145716
rect 253480 145528 253532 145580
rect 307116 145528 307168 145580
rect 184204 144984 184256 145036
rect 213920 144984 213972 145036
rect 303068 144984 303120 145036
rect 307484 144984 307536 145036
rect 174636 144916 174688 144968
rect 214012 144916 214064 144968
rect 279608 144916 279660 144968
rect 307668 144916 307720 144968
rect 252376 144848 252428 144900
rect 267832 144848 267884 144900
rect 324412 144848 324464 144900
rect 338212 144848 338264 144900
rect 252468 144780 252520 144832
rect 262496 144780 262548 144832
rect 324320 144780 324372 144832
rect 336740 144780 336792 144832
rect 290740 144236 290792 144288
rect 307576 144236 307628 144288
rect 253388 144168 253440 144220
rect 307392 144168 307444 144220
rect 304540 143624 304592 143676
rect 307668 143624 307720 143676
rect 167736 143556 167788 143608
rect 213920 143556 213972 143608
rect 257436 143556 257488 143608
rect 306564 143556 306616 143608
rect 252376 143488 252428 143540
rect 264980 143488 265032 143540
rect 324412 143488 324464 143540
rect 345020 143488 345072 143540
rect 252468 143420 252520 143472
rect 263692 143420 263744 143472
rect 324320 143420 324372 143472
rect 343824 143420 343876 143472
rect 251640 143352 251692 143404
rect 255320 143352 255372 143404
rect 322204 142332 322256 142384
rect 324412 142332 324464 142384
rect 202236 142196 202288 142248
rect 213920 142196 213972 142248
rect 276756 142196 276808 142248
rect 307668 142196 307720 142248
rect 173256 142128 173308 142180
rect 214012 142128 214064 142180
rect 253296 142128 253348 142180
rect 307576 142128 307628 142180
rect 324964 142128 325016 142180
rect 325700 142128 325752 142180
rect 252376 142060 252428 142112
rect 271972 142060 272024 142112
rect 324504 142060 324556 142112
rect 352012 142060 352064 142112
rect 324320 141992 324372 142044
rect 346492 141992 346544 142044
rect 294880 141380 294932 141432
rect 306472 141380 306524 141432
rect 252468 141108 252520 141160
rect 259552 141108 259604 141160
rect 210516 140836 210568 140888
rect 214012 140836 214064 140888
rect 171784 140768 171836 140820
rect 213920 140768 213972 140820
rect 251916 140768 251968 140820
rect 254860 140768 254912 140820
rect 252468 140700 252520 140752
rect 281724 140700 281776 140752
rect 324320 140700 324372 140752
rect 328736 140700 328788 140752
rect 252376 140632 252428 140684
rect 256976 140632 257028 140684
rect 180340 140020 180392 140072
rect 214564 140020 214616 140072
rect 252100 140020 252152 140072
rect 290464 140020 290516 140072
rect 282276 139476 282328 139528
rect 307300 139476 307352 139528
rect 207664 139408 207716 139460
rect 213920 139408 213972 139460
rect 267188 139408 267240 139460
rect 307668 139408 307720 139460
rect 252376 139340 252428 139392
rect 274732 139340 274784 139392
rect 324320 139340 324372 139392
rect 343732 139340 343784 139392
rect 252468 139272 252520 139324
rect 262312 139272 262364 139324
rect 324504 139272 324556 139324
rect 341064 139272 341116 139324
rect 294604 138116 294656 138168
rect 307300 138116 307352 138168
rect 278136 138048 278188 138100
rect 307668 138048 307720 138100
rect 196716 137980 196768 138032
rect 213920 137980 213972 138032
rect 250444 137980 250496 138032
rect 307576 137980 307628 138032
rect 252468 137912 252520 137964
rect 276112 137912 276164 137964
rect 324504 137912 324556 137964
rect 335636 137912 335688 137964
rect 252376 137844 252428 137896
rect 273444 137844 273496 137896
rect 324320 137844 324372 137896
rect 334164 137844 334216 137896
rect 177580 137232 177632 137284
rect 214564 137232 214616 137284
rect 254860 137232 254912 137284
rect 307024 137232 307076 137284
rect 2780 136960 2832 137012
rect 4804 136960 4856 137012
rect 292028 136688 292080 136740
rect 307576 136688 307628 136740
rect 166264 136620 166316 136672
rect 213920 136620 213972 136672
rect 250536 136620 250588 136672
rect 307668 136620 307720 136672
rect 252284 136552 252336 136604
rect 291936 136552 291988 136604
rect 324504 136552 324556 136604
rect 342260 136552 342312 136604
rect 252468 136484 252520 136536
rect 289176 136484 289228 136536
rect 252376 136416 252428 136468
rect 269764 136416 269816 136468
rect 252008 136348 252060 136400
rect 254584 136348 254636 136400
rect 324320 136348 324372 136400
rect 327264 136348 327316 136400
rect 300216 135464 300268 135516
rect 306748 135464 306800 135516
rect 289268 135396 289320 135448
rect 307668 135396 307720 135448
rect 285036 135328 285088 135380
rect 307484 135328 307536 135380
rect 178776 135260 178828 135312
rect 213920 135260 213972 135312
rect 265716 135260 265768 135312
rect 307576 135260 307628 135312
rect 252376 135192 252428 135244
rect 295984 135192 296036 135244
rect 324320 135192 324372 135244
rect 331404 135192 331456 135244
rect 252468 135124 252520 135176
rect 289084 135124 289136 135176
rect 286692 134512 286744 134564
rect 307392 134512 307444 134564
rect 181444 133900 181496 133952
rect 213920 133900 213972 133952
rect 293224 133900 293276 133952
rect 307668 133900 307720 133952
rect 252376 133832 252428 133884
rect 296076 133832 296128 133884
rect 324320 133832 324372 133884
rect 345204 133832 345256 133884
rect 252284 133764 252336 133816
rect 268384 133764 268436 133816
rect 252468 133696 252520 133748
rect 267004 133696 267056 133748
rect 295984 132608 296036 132660
rect 306564 132608 306616 132660
rect 202328 132540 202380 132592
rect 214012 132540 214064 132592
rect 287796 132540 287848 132592
rect 307116 132540 307168 132592
rect 173348 132472 173400 132524
rect 213920 132472 213972 132524
rect 273904 132472 273956 132524
rect 307668 132472 307720 132524
rect 252284 132404 252336 132456
rect 300124 132404 300176 132456
rect 252376 132336 252428 132388
rect 286416 132336 286468 132388
rect 252468 132268 252520 132320
rect 264428 132268 264480 132320
rect 203616 131180 203668 131232
rect 214012 131180 214064 131232
rect 286508 131180 286560 131232
rect 306932 131180 306984 131232
rect 171876 131112 171928 131164
rect 213920 131112 213972 131164
rect 283564 131112 283616 131164
rect 306564 131112 306616 131164
rect 252468 131044 252520 131096
rect 275376 131044 275428 131096
rect 324320 131044 324372 131096
rect 347872 131044 347924 131096
rect 252376 130976 252428 131028
rect 269856 130976 269908 131028
rect 324412 130976 324464 131028
rect 330024 130976 330076 131028
rect 252284 130908 252336 130960
rect 262864 130908 262916 130960
rect 269948 130364 270000 130416
rect 307300 130364 307352 130416
rect 290648 129820 290700 129872
rect 307484 129820 307536 129872
rect 171968 129752 172020 129804
rect 213920 129752 213972 129804
rect 275284 129752 275336 129804
rect 307668 129752 307720 129804
rect 252376 129684 252428 129736
rect 276664 129684 276716 129736
rect 324320 129684 324372 129736
rect 329932 129684 329984 129736
rect 252468 129616 252520 129668
rect 271328 129616 271380 129668
rect 324412 129616 324464 129668
rect 329840 129616 329892 129668
rect 290556 128460 290608 128512
rect 307484 128460 307536 128512
rect 280896 128392 280948 128444
rect 307576 128392 307628 128444
rect 176016 128324 176068 128376
rect 213920 128324 213972 128376
rect 252192 128324 252244 128376
rect 260196 128324 260248 128376
rect 271144 128324 271196 128376
rect 307668 128324 307720 128376
rect 252468 128256 252520 128308
rect 283748 128256 283800 128308
rect 324320 128256 324372 128308
rect 328552 128256 328604 128308
rect 252284 128188 252336 128240
rect 281080 128188 281132 128240
rect 252376 128120 252428 128172
rect 278228 128120 278280 128172
rect 283656 127100 283708 127152
rect 307576 127100 307628 127152
rect 282184 127032 282236 127084
rect 307668 127032 307720 127084
rect 198096 126964 198148 127016
rect 213920 126964 213972 127016
rect 280988 126964 281040 127016
rect 307484 126964 307536 127016
rect 252468 126896 252520 126948
rect 302884 126896 302936 126948
rect 251732 126828 251784 126880
rect 254860 126828 254912 126880
rect 252284 126216 252336 126268
rect 305736 126216 305788 126268
rect 207756 125672 207808 125724
rect 213920 125672 213972 125724
rect 289360 125672 289412 125724
rect 306564 125672 306616 125724
rect 59268 125604 59320 125656
rect 65156 125604 65208 125656
rect 176108 125604 176160 125656
rect 214012 125604 214064 125656
rect 254584 125604 254636 125656
rect 307668 125604 307720 125656
rect 252468 125536 252520 125588
rect 298836 125536 298888 125588
rect 324320 125536 324372 125588
rect 332692 125536 332744 125588
rect 252376 125468 252428 125520
rect 287980 125468 288032 125520
rect 302884 124380 302936 124432
rect 307668 124380 307720 124432
rect 298744 124312 298796 124364
rect 306564 124312 306616 124364
rect 187148 124244 187200 124296
rect 213920 124244 213972 124296
rect 287888 124244 287940 124296
rect 307484 124244 307536 124296
rect 62028 124176 62080 124228
rect 65524 124176 65576 124228
rect 169208 124176 169260 124228
rect 214012 124176 214064 124228
rect 255964 124176 256016 124228
rect 307576 124176 307628 124228
rect 252468 124108 252520 124160
rect 301504 124108 301556 124160
rect 324320 124108 324372 124160
rect 340972 124108 341024 124160
rect 252376 124040 252428 124092
rect 271236 124040 271288 124092
rect 324412 124040 324464 124092
rect 338396 124040 338448 124092
rect 252284 123972 252336 124024
rect 257528 123972 257580 124024
rect 301688 122952 301740 123004
rect 307668 122952 307720 123004
rect 170588 122884 170640 122936
rect 213920 122884 213972 122936
rect 289084 122884 289136 122936
rect 307484 122884 307536 122936
rect 61936 122816 61988 122868
rect 66076 122816 66128 122868
rect 169116 122816 169168 122868
rect 214012 122816 214064 122868
rect 272524 122816 272576 122868
rect 307576 122816 307628 122868
rect 252468 122748 252520 122800
rect 297456 122748 297508 122800
rect 324320 122748 324372 122800
rect 358820 122748 358872 122800
rect 252284 122680 252336 122732
rect 264244 122680 264296 122732
rect 252376 122408 252428 122460
rect 258908 122408 258960 122460
rect 297364 121592 297416 121644
rect 307484 121592 307536 121644
rect 209228 121524 209280 121576
rect 214012 121524 214064 121576
rect 293316 121524 293368 121576
rect 307576 121524 307628 121576
rect 177396 121456 177448 121508
rect 213920 121456 213972 121508
rect 267004 121456 267056 121508
rect 307668 121456 307720 121508
rect 252376 121388 252428 121440
rect 291844 121388 291896 121440
rect 324320 121388 324372 121440
rect 356060 121388 356112 121440
rect 252468 121320 252520 121372
rect 265624 121320 265676 121372
rect 252468 120912 252520 120964
rect 258724 120912 258776 120964
rect 296076 120232 296128 120284
rect 307668 120232 307720 120284
rect 188436 120164 188488 120216
rect 213920 120164 213972 120216
rect 286416 120164 286468 120216
rect 307576 120164 307628 120216
rect 166356 120096 166408 120148
rect 214012 120096 214064 120148
rect 271236 120096 271288 120148
rect 307116 120096 307168 120148
rect 252468 120028 252520 120080
rect 262956 120028 263008 120080
rect 252284 119960 252336 120012
rect 253480 119960 253532 120012
rect 252376 119348 252428 119400
rect 293408 119348 293460 119400
rect 170404 118804 170456 118856
rect 213920 118804 213972 118856
rect 304264 118804 304316 118856
rect 307668 118804 307720 118856
rect 185676 118736 185728 118788
rect 214012 118736 214064 118788
rect 291844 118736 291896 118788
rect 307576 118736 307628 118788
rect 262864 118668 262916 118720
rect 307116 118668 307168 118720
rect 252468 118600 252520 118652
rect 264336 118600 264388 118652
rect 324412 118600 324464 118652
rect 345112 118600 345164 118652
rect 324320 118532 324372 118584
rect 339684 118532 339736 118584
rect 252468 117648 252520 117700
rect 258816 117648 258868 117700
rect 300124 117512 300176 117564
rect 306564 117512 306616 117564
rect 298836 117444 298888 117496
rect 307668 117444 307720 117496
rect 174728 117376 174780 117428
rect 214012 117376 214064 117428
rect 265624 117376 265676 117428
rect 307576 117376 307628 117428
rect 170680 117308 170732 117360
rect 213920 117308 213972 117360
rect 264244 117308 264296 117360
rect 307116 117308 307168 117360
rect 252468 117240 252520 117292
rect 282460 117240 282512 117292
rect 324320 117240 324372 117292
rect 338304 117240 338356 117292
rect 252376 117172 252428 117224
rect 268476 117172 268528 117224
rect 296352 116560 296404 116612
rect 307024 116560 307076 116612
rect 252468 116492 252520 116544
rect 260104 116492 260156 116544
rect 198188 116016 198240 116068
rect 214012 116016 214064 116068
rect 282368 116016 282420 116068
rect 306932 116016 306984 116068
rect 181536 115948 181588 116000
rect 213920 115948 213972 116000
rect 268384 115948 268436 116000
rect 307668 115948 307720 116000
rect 252376 115880 252428 115932
rect 267096 115880 267148 115932
rect 324412 115880 324464 115932
rect 351920 115880 351972 115932
rect 324320 115812 324372 115864
rect 342444 115812 342496 115864
rect 169024 115268 169076 115320
rect 203524 115268 203576 115320
rect 173440 115200 173492 115252
rect 214656 115200 214708 115252
rect 252468 115200 252520 115252
rect 297640 115200 297692 115252
rect 297548 114656 297600 114708
rect 307668 114656 307720 114708
rect 294696 114588 294748 114640
rect 307576 114588 307628 114640
rect 211896 114520 211948 114572
rect 213920 114520 213972 114572
rect 269764 114520 269816 114572
rect 307116 114520 307168 114572
rect 252468 114452 252520 114504
rect 275468 114452 275520 114504
rect 324412 114452 324464 114504
rect 335452 114452 335504 114504
rect 252284 114384 252336 114436
rect 256148 114384 256200 114436
rect 324320 114384 324372 114436
rect 333980 114384 334032 114436
rect 251732 114316 251784 114368
rect 254768 114316 254820 114368
rect 284944 113296 284996 113348
rect 307576 113296 307628 113348
rect 276664 113228 276716 113280
rect 307668 113228 307720 113280
rect 180248 113160 180300 113212
rect 213920 113160 213972 113212
rect 260104 113160 260156 113212
rect 307484 113160 307536 113212
rect 252468 113092 252520 113144
rect 300400 113092 300452 113144
rect 324320 113092 324372 113144
rect 339500 113092 339552 113144
rect 252100 112412 252152 112464
rect 303068 112412 303120 112464
rect 252468 112276 252520 112328
rect 259000 112276 259052 112328
rect 301504 111936 301556 111988
rect 307668 111936 307720 111988
rect 189816 111868 189868 111920
rect 214012 111868 214064 111920
rect 302976 111868 303028 111920
rect 307576 111868 307628 111920
rect 170496 111800 170548 111852
rect 213920 111800 213972 111852
rect 297456 111800 297508 111852
rect 307668 111800 307720 111852
rect 3148 111732 3200 111784
rect 11704 111732 11756 111784
rect 168288 111732 168340 111784
rect 199568 111732 199620 111784
rect 252468 111732 252520 111784
rect 296168 111732 296220 111784
rect 324320 111732 324372 111784
rect 340880 111732 340932 111784
rect 252376 111664 252428 111716
rect 272800 111664 272852 111716
rect 304448 110576 304500 110628
rect 307484 110576 307536 110628
rect 177488 110508 177540 110560
rect 213920 110508 213972 110560
rect 252192 110508 252244 110560
rect 256240 110508 256292 110560
rect 296260 110508 296312 110560
rect 307668 110508 307720 110560
rect 166448 110440 166500 110492
rect 214012 110440 214064 110492
rect 272708 110440 272760 110492
rect 307576 110440 307628 110492
rect 167828 110372 167880 110424
rect 177580 110372 177632 110424
rect 252376 110372 252428 110424
rect 300308 110372 300360 110424
rect 324412 110372 324464 110424
rect 336832 110372 336884 110424
rect 252468 110304 252520 110356
rect 273996 110304 274048 110356
rect 324320 110304 324372 110356
rect 332600 110304 332652 110356
rect 252284 110236 252336 110288
rect 256056 110236 256108 110288
rect 301596 109148 301648 109200
rect 307484 109148 307536 109200
rect 195520 109080 195572 109132
rect 214012 109080 214064 109132
rect 298928 109080 298980 109132
rect 307576 109080 307628 109132
rect 169024 109012 169076 109064
rect 213920 109012 213972 109064
rect 275376 109012 275428 109064
rect 307668 109012 307720 109064
rect 168104 108944 168156 108996
rect 180340 108944 180392 108996
rect 252376 108944 252428 108996
rect 301780 108944 301832 108996
rect 324320 108944 324372 108996
rect 342536 108944 342588 108996
rect 252468 108876 252520 108928
rect 297732 108876 297784 108928
rect 251732 108808 251784 108860
rect 254676 108808 254728 108860
rect 178960 108264 179012 108316
rect 214748 108264 214800 108316
rect 297640 107856 297692 107908
rect 307668 107856 307720 107908
rect 300400 107720 300452 107772
rect 307484 107720 307536 107772
rect 182916 107652 182968 107704
rect 213920 107652 213972 107704
rect 303068 107652 303120 107704
rect 307576 107652 307628 107704
rect 252376 107584 252428 107636
rect 305644 107584 305696 107636
rect 252468 107516 252520 107568
rect 304356 107516 304408 107568
rect 252284 107448 252336 107500
rect 257344 107448 257396 107500
rect 177580 106360 177632 106412
rect 213920 106360 213972 106412
rect 301780 106360 301832 106412
rect 307668 106360 307720 106412
rect 167828 106292 167880 106344
rect 214012 106292 214064 106344
rect 304632 106292 304684 106344
rect 306748 106292 306800 106344
rect 252468 106224 252520 106276
rect 261484 106224 261536 106276
rect 324320 106224 324372 106276
rect 352104 106224 352156 106276
rect 251180 106156 251232 106208
rect 253388 106156 253440 106208
rect 252376 105476 252428 105528
rect 304540 105544 304592 105596
rect 258724 105000 258776 105052
rect 307668 105000 307720 105052
rect 188528 104864 188580 104916
rect 213920 104864 213972 104916
rect 303160 104864 303212 104916
rect 307576 104864 307628 104916
rect 252468 104796 252520 104848
rect 290740 104796 290792 104848
rect 173164 104116 173216 104168
rect 216220 104116 216272 104168
rect 279608 104116 279660 104168
rect 252468 103980 252520 104032
rect 304356 103640 304408 103692
rect 307484 103640 307536 103692
rect 206560 103572 206612 103624
rect 214012 103572 214064 103624
rect 290464 103572 290516 103624
rect 307576 103572 307628 103624
rect 192576 103504 192628 103556
rect 213920 103504 213972 103556
rect 279516 103504 279568 103556
rect 307668 103504 307720 103556
rect 324504 103436 324556 103488
rect 357440 103436 357492 103488
rect 324320 103300 324372 103352
rect 324688 103300 324740 103352
rect 252284 103164 252336 103216
rect 253296 103164 253348 103216
rect 324320 103164 324372 103216
rect 327080 103164 327132 103216
rect 252192 103096 252244 103148
rect 257436 103096 257488 103148
rect 289176 102280 289228 102332
rect 307576 102280 307628 102332
rect 203708 102212 203760 102264
rect 213920 102212 213972 102264
rect 257344 102212 257396 102264
rect 307668 102212 307720 102264
rect 199568 102144 199620 102196
rect 214012 102144 214064 102196
rect 253388 102144 253440 102196
rect 307484 102144 307536 102196
rect 252468 102076 252520 102128
rect 276756 102076 276808 102128
rect 169300 101396 169352 101448
rect 214472 101396 214524 101448
rect 252192 101396 252244 101448
rect 267188 101396 267240 101448
rect 267096 100920 267148 100972
rect 307576 100920 307628 100972
rect 293408 100852 293460 100904
rect 307668 100852 307720 100904
rect 206468 100784 206520 100836
rect 214012 100784 214064 100836
rect 273996 100784 274048 100836
rect 307484 100784 307536 100836
rect 173164 100716 173216 100768
rect 213920 100716 213972 100768
rect 252284 100648 252336 100700
rect 296352 100648 296404 100700
rect 324320 100648 324372 100700
rect 331496 100648 331548 100700
rect 468484 100648 468536 100700
rect 580172 100648 580224 100700
rect 252468 100580 252520 100632
rect 294880 100580 294932 100632
rect 252376 100512 252428 100564
rect 269948 100512 270000 100564
rect 300308 99492 300360 99544
rect 306748 99492 306800 99544
rect 296168 99424 296220 99476
rect 307668 99424 307720 99476
rect 294788 99356 294840 99408
rect 307576 99356 307628 99408
rect 252468 99220 252520 99272
rect 264520 99220 264572 99272
rect 252376 99152 252428 99204
rect 286692 99152 286744 99204
rect 166540 98064 166592 98116
rect 214012 98064 214064 98116
rect 286600 98064 286652 98116
rect 307576 98064 307628 98116
rect 164884 97996 164936 98048
rect 213920 97996 213972 98048
rect 261484 97996 261536 98048
rect 307668 97996 307720 98048
rect 3516 97928 3568 97980
rect 17224 97928 17276 97980
rect 167920 97248 167972 97300
rect 214104 97248 214156 97300
rect 252468 97248 252520 97300
rect 272616 97248 272668 97300
rect 291936 96772 291988 96824
rect 307668 96772 307720 96824
rect 278228 96704 278280 96756
rect 306932 96704 306984 96756
rect 253204 96636 253256 96688
rect 307668 96636 307720 96688
rect 199476 96568 199528 96620
rect 321284 96568 321336 96620
rect 286324 96500 286376 96552
rect 321468 96500 321520 96552
rect 249064 95208 249116 95260
rect 306932 95208 306984 95260
rect 210424 95140 210476 95192
rect 324412 95140 324464 95192
rect 216128 95072 216180 95124
rect 324688 95072 324740 95124
rect 59268 95004 59320 95056
rect 206560 95004 206612 95056
rect 308496 95004 308548 95056
rect 321560 95004 321612 95056
rect 162860 94528 162912 94580
rect 203616 94528 203668 94580
rect 122840 94460 122892 94512
rect 214656 94460 214708 94512
rect 151728 93916 151780 93968
rect 178868 93916 178920 93968
rect 129372 93848 129424 93900
rect 167736 93848 167788 93900
rect 151728 93440 151780 93492
rect 175924 93440 175976 93492
rect 135720 93372 135772 93424
rect 167644 93372 167696 93424
rect 120632 93304 120684 93356
rect 170588 93304 170640 93356
rect 115480 93236 115532 93288
rect 166264 93236 166316 93288
rect 85672 93168 85724 93220
rect 164884 93168 164936 93220
rect 126612 93100 126664 93152
rect 214840 93100 214892 93152
rect 238024 93100 238076 93152
rect 251180 93100 251232 93152
rect 74816 92420 74868 92472
rect 214748 92420 214800 92472
rect 88984 92352 89036 92404
rect 167920 92352 167972 92404
rect 95056 92284 95108 92336
rect 122840 92284 122892 92336
rect 134432 92284 134484 92336
rect 210608 92284 210660 92336
rect 105544 92216 105596 92268
rect 126612 92216 126664 92268
rect 126704 92216 126756 92268
rect 202236 92216 202288 92268
rect 116768 92148 116820 92200
rect 169300 92148 169352 92200
rect 128176 92080 128228 92132
rect 173440 92080 173492 92132
rect 178684 91740 178736 91792
rect 307300 91740 307352 91792
rect 102048 91060 102100 91112
rect 118700 91060 118752 91112
rect 67364 90992 67416 91044
rect 203708 90992 203760 91044
rect 62028 90924 62080 90976
rect 192576 90924 192628 90976
rect 106648 90856 106700 90908
rect 173348 90856 173400 90908
rect 110328 90788 110380 90840
rect 170680 90788 170732 90840
rect 124036 90720 124088 90772
rect 169208 90720 169260 90772
rect 151728 90652 151780 90704
rect 177304 90652 177356 90704
rect 115572 89632 115624 89684
rect 213368 89632 213420 89684
rect 113824 89564 113876 89616
rect 185676 89564 185728 89616
rect 118700 89496 118752 89548
rect 189816 89496 189868 89548
rect 126888 89428 126940 89480
rect 176108 89428 176160 89480
rect 125416 89360 125468 89412
rect 171784 89360 171836 89412
rect 153016 89292 153068 89344
rect 184296 89292 184348 89344
rect 188344 88952 188396 89004
rect 324320 88952 324372 89004
rect 107200 88272 107252 88324
rect 211896 88272 211948 88324
rect 90732 88204 90784 88256
rect 188528 88204 188580 88256
rect 100208 88136 100260 88188
rect 166448 88136 166500 88188
rect 118240 88068 118292 88120
rect 177396 88068 177448 88120
rect 132408 88000 132460 88052
rect 174636 88000 174688 88052
rect 188344 87592 188396 87644
rect 307208 87592 307260 87644
rect 67640 86912 67692 86964
rect 214564 86912 214616 86964
rect 97080 86844 97132 86896
rect 198096 86844 198148 86896
rect 108488 86776 108540 86828
rect 181536 86776 181588 86828
rect 117136 86708 117188 86760
rect 166356 86708 166408 86760
rect 126704 86640 126756 86692
rect 173256 86640 173308 86692
rect 202144 86232 202196 86284
rect 307760 86232 307812 86284
rect 3516 85484 3568 85536
rect 54484 85484 54536 85536
rect 102968 85484 103020 85536
rect 213460 85484 213512 85536
rect 108212 85416 108264 85468
rect 202328 85416 202380 85468
rect 109592 85348 109644 85400
rect 181444 85348 181496 85400
rect 122840 85280 122892 85332
rect 187148 85280 187200 85332
rect 112536 85212 112588 85264
rect 170404 85212 170456 85264
rect 133236 85144 133288 85196
rect 174544 85144 174596 85196
rect 206284 84804 206336 84856
rect 324412 84804 324464 84856
rect 67548 84124 67600 84176
rect 206468 84124 206520 84176
rect 115848 84056 115900 84108
rect 188436 84056 188488 84108
rect 96528 83988 96580 84040
rect 169024 83988 169076 84040
rect 111708 83920 111760 83972
rect 174728 83920 174780 83972
rect 196624 83444 196676 83496
rect 314660 83444 314712 83496
rect 110144 82764 110196 82816
rect 198188 82764 198240 82816
rect 124128 82696 124180 82748
rect 210516 82696 210568 82748
rect 99196 82628 99248 82680
rect 177488 82628 177540 82680
rect 101956 82560 102008 82612
rect 171968 82560 172020 82612
rect 122656 82492 122708 82544
rect 169116 82492 169168 82544
rect 206376 82084 206428 82136
rect 329840 82084 329892 82136
rect 92388 81336 92440 81388
rect 177580 81336 177632 81388
rect 125508 81268 125560 81320
rect 207756 81268 207808 81320
rect 100668 81200 100720 81252
rect 170496 81200 170548 81252
rect 104716 81132 104768 81184
rect 171876 81132 171928 81184
rect 131028 81064 131080 81116
rect 184204 81064 184256 81116
rect 209044 80656 209096 80708
rect 325700 80656 325752 80708
rect 119988 79976 120040 80028
rect 209228 79976 209280 80028
rect 95148 79908 95200 79960
rect 182916 79908 182968 79960
rect 86868 79840 86920 79892
rect 166540 79840 166592 79892
rect 118608 79772 118660 79824
rect 196716 79772 196768 79824
rect 97908 78616 97960 78668
rect 195520 78616 195572 78668
rect 122748 78548 122800 78600
rect 213276 78548 213328 78600
rect 93768 78480 93820 78532
rect 167828 78480 167880 78532
rect 101864 78412 101916 78464
rect 176016 78412 176068 78464
rect 211804 78004 211856 78056
rect 260840 78004 260892 78056
rect 280804 78004 280856 78056
rect 316040 78004 316092 78056
rect 180064 77936 180116 77988
rect 321560 77936 321612 77988
rect 85488 77188 85540 77240
rect 173164 77188 173216 77240
rect 121368 77120 121420 77172
rect 207664 77120 207716 77172
rect 114468 77052 114520 77104
rect 178776 77052 178828 77104
rect 92480 76508 92532 76560
rect 300216 76508 300268 76560
rect 104808 75828 104860 75880
rect 180248 75828 180300 75880
rect 95240 75216 95292 75268
rect 265716 75216 265768 75268
rect 69020 75148 69072 75200
rect 303160 75148 303212 75200
rect 122840 73924 122892 73976
rect 254584 73924 254636 73976
rect 99380 73856 99432 73908
rect 285036 73856 285088 73908
rect 71780 73788 71832 73840
rect 305920 73788 305972 73840
rect 115940 72564 115992 72616
rect 255964 72564 256016 72616
rect 84200 72496 84252 72548
rect 271236 72496 271288 72548
rect 67640 72428 67692 72480
rect 273904 72428 273956 72480
rect 98000 71068 98052 71120
rect 301688 71068 301740 71120
rect 46940 71000 46992 71052
rect 253388 71000 253440 71052
rect 110420 69708 110472 69760
rect 292028 69708 292080 69760
rect 75920 69640 75972 69692
rect 304632 69640 304684 69692
rect 113180 68416 113232 68468
rect 294604 68416 294656 68468
rect 78680 68348 78732 68400
rect 301780 68348 301832 68400
rect 4160 68280 4212 68332
rect 249064 68280 249116 68332
rect 82820 66920 82872 66972
rect 300400 66920 300452 66972
rect 13820 66852 13872 66904
rect 289360 66852 289412 66904
rect 85580 65560 85632 65612
rect 305828 65560 305880 65612
rect 60740 65492 60792 65544
rect 286508 65492 286560 65544
rect 89720 64132 89772 64184
rect 303068 64132 303120 64184
rect 93860 62772 93912 62824
rect 297640 62772 297692 62824
rect 96620 61412 96672 61464
rect 275376 61412 275428 61464
rect 278044 61412 278096 61464
rect 316132 61412 316184 61464
rect 44180 61344 44232 61396
rect 282368 61344 282420 61396
rect 185584 60052 185636 60104
rect 313280 60052 313332 60104
rect 12440 59984 12492 60036
rect 276664 59984 276716 60036
rect 3056 59304 3108 59356
rect 53104 59304 53156 59356
rect 100760 58692 100812 58744
rect 298928 58692 298980 58744
rect 52460 58624 52512 58676
rect 290648 58624 290700 58676
rect 103520 57264 103572 57316
rect 301596 57264 301648 57316
rect 37280 57196 37332 57248
rect 269764 57196 269816 57248
rect 107660 55904 107712 55956
rect 296260 55904 296312 55956
rect 34520 55836 34572 55888
rect 294696 55836 294748 55888
rect 110512 54544 110564 54596
rect 304448 54544 304500 54596
rect 30380 54476 30432 54528
rect 297548 54476 297600 54528
rect 114560 53048 114612 53100
rect 272708 53048 272760 53100
rect 124220 51756 124272 51808
rect 282276 51756 282328 51808
rect 16580 51688 16632 51740
rect 300308 51688 300360 51740
rect 81440 50396 81492 50448
rect 293224 50396 293276 50448
rect 27620 50328 27672 50380
rect 260104 50328 260156 50380
rect 106280 49104 106332 49156
rect 250536 49104 250588 49156
rect 121460 49036 121512 49088
rect 302976 49036 303028 49088
rect 17960 48968 18012 49020
rect 284944 48968 284996 49020
rect 31760 47608 31812 47660
rect 290556 47608 290608 47660
rect 20720 47540 20772 47592
rect 294788 47540 294840 47592
rect 180156 46860 180208 46912
rect 580172 46860 580224 46912
rect 73160 46248 73212 46300
rect 262864 46248 262916 46300
rect 93952 46180 94004 46232
rect 293316 46180 293368 46232
rect 3424 45500 3476 45552
rect 15844 45500 15896 45552
rect 35900 44888 35952 44940
rect 271144 44888 271196 44940
rect 26240 44820 26292 44872
rect 293408 44820 293460 44872
rect 88340 43460 88392 43512
rect 289268 43460 289320 43512
rect 29000 43392 29052 43444
rect 273996 43392 274048 43444
rect 27712 42100 27764 42152
rect 280988 42100 281040 42152
rect 33140 42032 33192 42084
rect 305736 42032 305788 42084
rect 38660 40740 38712 40792
rect 280896 40740 280948 40792
rect 11060 40672 11112 40724
rect 296168 40672 296220 40724
rect 51080 39380 51132 39432
rect 279516 39380 279568 39432
rect 23480 39312 23532 39364
rect 283656 39312 283708 39364
rect 45560 37952 45612 38004
rect 275284 37952 275336 38004
rect 6920 37884 6972 37936
rect 286600 37884 286652 37936
rect 11152 36524 11204 36576
rect 278228 36524 278280 36576
rect 57888 35844 57940 35896
rect 251180 35844 251232 35896
rect 109040 35232 109092 35284
rect 287888 35232 287940 35284
rect 4804 35164 4856 35216
rect 57888 35164 57940 35216
rect 85672 35164 85724 35216
rect 308588 35164 308640 35216
rect 1308 34416 1360 34468
rect 249156 34416 249208 34468
rect 63500 33736 63552 33788
rect 283564 33736 283616 33788
rect 20 33124 72 33176
rect 1308 33124 1360 33176
rect 3516 33056 3568 33108
rect 43444 33056 43496 33108
rect 77300 32444 77352 32496
rect 296076 32444 296128 32496
rect 37188 32376 37240 32428
rect 270500 32376 270552 32428
rect 70400 31016 70452 31068
rect 287796 31016 287848 31068
rect 195244 29724 195296 29776
rect 251180 29724 251232 29776
rect 2872 29656 2924 29708
rect 253204 29656 253256 29708
rect 43444 29588 43496 29640
rect 307116 29588 307168 29640
rect 182824 28296 182876 28348
rect 262220 28296 262272 28348
rect 8300 28228 8352 28280
rect 301504 28228 301556 28280
rect 118700 26936 118752 26988
rect 297456 26936 297508 26988
rect 59360 26868 59412 26920
rect 265624 26868 265676 26920
rect 120080 25644 120132 25696
rect 250444 25644 250496 25696
rect 86960 25576 87012 25628
rect 297364 25576 297416 25628
rect 57980 25508 58032 25560
rect 304356 25508 304408 25560
rect 204996 24216 205048 24268
rect 244280 24216 244332 24268
rect 193864 24148 193916 24200
rect 292580 24148 292632 24200
rect 102140 24080 102192 24132
rect 272524 24080 272576 24132
rect 69112 22788 69164 22840
rect 291844 22788 291896 22840
rect 19340 22720 19392 22772
rect 261484 22720 261536 22772
rect 189724 21496 189776 21548
rect 309140 21496 309192 21548
rect 62120 21428 62172 21480
rect 300124 21428 300176 21480
rect 34428 21360 34480 21412
rect 280160 21360 280212 21412
rect 3424 20612 3476 20664
rect 40684 20612 40736 20664
rect 91100 19932 91152 19984
rect 267004 19932 267056 19984
rect 191104 18708 191156 18760
rect 241520 18708 241572 18760
rect 35992 18640 36044 18692
rect 267096 18640 267148 18692
rect 55220 18572 55272 18624
rect 298836 18572 298888 18624
rect 64788 17348 64840 17400
rect 242992 17348 243044 17400
rect 111800 17280 111852 17332
rect 302884 17280 302936 17332
rect 74540 17212 74592 17264
rect 295984 17212 296036 17264
rect 195428 15988 195480 16040
rect 295616 15988 295668 16040
rect 209136 15920 209188 15972
rect 322940 15920 322992 15972
rect 48504 15852 48556 15904
rect 268384 15852 268436 15904
rect 192484 14560 192536 14612
rect 306380 14560 306432 14612
rect 40224 14492 40276 14544
rect 257344 14492 257396 14544
rect 54944 14424 54996 14476
rect 290464 14424 290516 14476
rect 216220 13132 216272 13184
rect 259460 13132 259512 13184
rect 203524 13064 203576 13116
rect 267740 13064 267792 13116
rect 187056 11840 187108 11892
rect 247592 11840 247644 11892
rect 191196 11772 191248 11824
rect 328000 11772 328052 11824
rect 80888 11704 80940 11756
rect 286416 11704 286468 11756
rect 186964 10412 187016 10464
rect 256700 10412 256752 10464
rect 52552 10344 52604 10396
rect 264244 10344 264296 10396
rect 44272 10276 44324 10328
rect 289176 10276 289228 10328
rect 200764 9052 200816 9104
rect 254676 9052 254728 9104
rect 119896 8984 119948 9036
rect 298744 8984 298796 9036
rect 41880 8916 41932 8968
rect 307024 8916 307076 8968
rect 216036 7692 216088 7744
rect 239312 7692 239364 7744
rect 39948 7624 40000 7676
rect 168380 7624 168432 7676
rect 198004 7624 198056 7676
rect 249984 7624 250036 7676
rect 4068 7556 4120 7608
rect 25504 7556 25556 7608
rect 105728 7556 105780 7608
rect 289084 7556 289136 7608
rect 199384 6264 199436 6316
rect 292580 6264 292632 6316
rect 65524 6196 65576 6248
rect 305644 6196 305696 6248
rect 19432 6128 19484 6180
rect 282184 6128 282236 6180
rect 117596 4836 117648 4888
rect 278136 4836 278188 4888
rect 62028 4768 62080 4820
rect 258724 4768 258776 4820
rect 309692 4088 309744 4140
rect 318524 4088 318576 4140
rect 217324 3612 217376 3664
rect 242900 3612 242952 3664
rect 308404 3612 308456 3664
rect 320916 3680 320968 3732
rect 316132 3612 316184 3664
rect 317328 3612 317380 3664
rect 1676 3544 1728 3596
rect 4804 3544 4856 3596
rect 125876 3544 125928 3596
rect 171140 3544 171192 3596
rect 213184 3544 213236 3596
rect 240508 3544 240560 3596
rect 251180 3544 251232 3596
rect 252376 3544 252428 3596
rect 259460 3544 259512 3596
rect 260656 3544 260708 3596
rect 299480 3544 299532 3596
rect 300768 3544 300820 3596
rect 307852 3544 307904 3596
rect 309048 3544 309100 3596
rect 309876 3544 309928 3596
rect 329196 3544 329248 3596
rect 11060 3476 11112 3528
rect 11980 3476 12032 3528
rect 25320 3476 25372 3528
rect 43444 3476 43496 3528
rect 44180 3476 44232 3528
rect 45100 3476 45152 3528
rect 52460 3476 52512 3528
rect 53380 3476 53432 3528
rect 85580 3476 85632 3528
rect 86500 3476 86552 3528
rect 103336 3476 103388 3528
rect 188344 3476 188396 3528
rect 215944 3476 215996 3528
rect 253480 3476 253532 3528
rect 287704 3476 287756 3528
rect 312636 3476 312688 3528
rect 324412 3476 324464 3528
rect 325608 3476 325660 3528
rect 349160 3476 349212 3528
rect 350448 3476 350500 3528
rect 6460 3408 6512 3460
rect 15200 3408 15252 3460
rect 43076 3408 43128 3460
rect 178684 3408 178736 3460
rect 204904 3408 204956 3460
rect 246396 3408 246448 3460
rect 279424 3408 279476 3460
rect 311440 3408 311492 3460
rect 342168 3408 342220 3460
rect 353300 3408 353352 3460
rect 235816 2932 235868 2984
rect 238024 2932 238076 2984
rect 66720 2116 66772 2168
rect 304264 2116 304316 2168
rect 15936 2048 15988 2100
rect 291936 2048 291988 2100
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 700262 8156 703520
rect 8116 700256 8168 700262
rect 8116 700198 8168 700204
rect 14464 700256 14516 700262
rect 14464 700198 14516 700204
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3422 632088 3478 632097
rect 3422 632023 3478 632032
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3238 566944 3294 566953
rect 3238 566879 3294 566888
rect 3252 565894 3280 566879
rect 3240 565888 3292 565894
rect 3240 565830 3292 565836
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2976 527202 3004 527847
rect 2964 527196 3016 527202
rect 2964 527138 3016 527144
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3054 475688 3110 475697
rect 3054 475623 3110 475632
rect 3068 474774 3096 475623
rect 3056 474768 3108 474774
rect 3056 474710 3108 474716
rect 2778 462632 2834 462641
rect 2778 462567 2780 462576
rect 2832 462567 2834 462576
rect 2780 462538 2832 462544
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 2870 410544 2926 410553
rect 2870 410479 2926 410488
rect 2884 409902 2912 410479
rect 2872 409896 2924 409902
rect 2872 409838 2924 409844
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3344 371278 3372 371311
rect 3332 371272 3384 371278
rect 3332 371214 3384 371220
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3344 357474 3372 358391
rect 3332 357468 3384 357474
rect 3332 357410 3384 357416
rect 3332 346384 3384 346390
rect 3332 346326 3384 346332
rect 3344 345409 3372 346326
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3436 334626 3464 632023
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618322 3556 619103
rect 3516 618316 3568 618322
rect 3516 618258 3568 618264
rect 3514 606112 3570 606121
rect 3514 606047 3570 606056
rect 3528 605878 3556 606047
rect 3516 605872 3568 605878
rect 3516 605814 3568 605820
rect 3514 553888 3570 553897
rect 3514 553823 3516 553832
rect 3568 553823 3570 553832
rect 7564 553852 7616 553858
rect 3516 553794 3568 553800
rect 7564 553794 7616 553800
rect 7576 530602 7604 553794
rect 7564 530596 7616 530602
rect 7564 530538 7616 530544
rect 7564 527196 7616 527202
rect 7564 527138 7616 527144
rect 3514 514856 3570 514865
rect 3514 514791 3516 514800
rect 3568 514791 3570 514800
rect 3516 514762 3568 514768
rect 4804 462596 4856 462602
rect 4804 462538 4856 462544
rect 3514 423600 3570 423609
rect 3514 423535 3570 423544
rect 3528 422346 3556 423535
rect 3516 422340 3568 422346
rect 3516 422282 3568 422288
rect 3516 397520 3568 397526
rect 3514 397488 3516 397497
rect 3568 397488 3570 397497
rect 3514 397423 3570 397432
rect 3516 374672 3568 374678
rect 3516 374614 3568 374620
rect 3424 334620 3476 334626
rect 3424 334562 3476 334568
rect 3528 319297 3556 374614
rect 4816 339454 4844 462538
rect 7576 391270 7604 527138
rect 11704 448588 11756 448594
rect 11704 448530 11756 448536
rect 7564 391264 7616 391270
rect 7564 391206 7616 391212
rect 4804 339448 4856 339454
rect 4804 339390 4856 339396
rect 3514 319288 3570 319297
rect 3514 319223 3570 319232
rect 3528 316034 3556 319223
rect 3436 316006 3556 316034
rect 3436 312594 3464 316006
rect 3424 312588 3476 312594
rect 3424 312530 3476 312536
rect 3424 306332 3476 306338
rect 3424 306274 3476 306280
rect 3436 306241 3464 306274
rect 3422 306232 3478 306241
rect 3422 306167 3478 306176
rect 3424 296812 3476 296818
rect 3424 296754 3476 296760
rect 3330 267200 3386 267209
rect 3330 267135 3332 267144
rect 3384 267135 3386 267144
rect 3332 267106 3384 267112
rect 3148 255264 3200 255270
rect 3148 255206 3200 255212
rect 3160 254153 3188 255206
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3054 241088 3110 241097
rect 3054 241023 3110 241032
rect 3068 240174 3096 241023
rect 3056 240168 3108 240174
rect 3056 240110 3108 240116
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 1306 200696 1362 200705
rect 1306 200631 1362 200640
rect 1320 34474 1348 200631
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 2780 137012 2832 137018
rect 2780 136954 2832 136960
rect 2792 136785 2820 136954
rect 2778 136776 2834 136785
rect 2778 136711 2834 136720
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3436 71641 3464 296754
rect 11716 296002 11744 448530
rect 14476 399498 14504 700198
rect 24320 698970 24348 703520
rect 24308 698964 24360 698970
rect 24308 698906 24360 698912
rect 35164 656940 35216 656946
rect 35164 656882 35216 656888
rect 15844 618316 15896 618322
rect 15844 618258 15896 618264
rect 15856 400926 15884 618258
rect 25504 605872 25556 605878
rect 25504 605814 25556 605820
rect 15844 400920 15896 400926
rect 15844 400862 15896 400868
rect 14464 399492 14516 399498
rect 14464 399434 14516 399440
rect 15200 397520 15252 397526
rect 15200 397462 15252 397468
rect 15212 396778 15240 397462
rect 15200 396772 15252 396778
rect 15200 396714 15252 396720
rect 21364 382288 21416 382294
rect 21364 382230 21416 382236
rect 21376 346390 21404 382230
rect 22744 357468 22796 357474
rect 22744 357410 22796 357416
rect 21364 346384 21416 346390
rect 21364 346326 21416 346332
rect 22756 344350 22784 357410
rect 22744 344344 22796 344350
rect 22744 344286 22796 344292
rect 25516 333878 25544 605814
rect 32404 579692 32456 579698
rect 32404 579634 32456 579640
rect 32416 338094 32444 579634
rect 35176 453354 35204 656882
rect 35256 474768 35308 474774
rect 35256 474710 35308 474716
rect 35164 453348 35216 453354
rect 35164 453290 35216 453296
rect 34336 379704 34388 379710
rect 34336 379646 34388 379652
rect 32404 338088 32456 338094
rect 32404 338030 32456 338036
rect 25504 333872 25556 333878
rect 25504 333814 25556 333820
rect 11704 295996 11756 296002
rect 11704 295938 11756 295944
rect 14464 294636 14516 294642
rect 14464 294578 14516 294584
rect 3608 293276 3660 293282
rect 3608 293218 3660 293224
rect 3514 293176 3570 293185
rect 3514 293111 3570 293120
rect 3528 292602 3556 293111
rect 3516 292596 3568 292602
rect 3516 292538 3568 292544
rect 3620 277394 3648 293218
rect 11704 292596 11756 292602
rect 11704 292538 11756 292544
rect 3528 277366 3648 277394
rect 3528 188873 3556 277366
rect 7564 267164 7616 267170
rect 7564 267106 7616 267112
rect 4804 257372 4856 257378
rect 4804 257314 4856 257320
rect 3608 225616 3660 225622
rect 3608 225558 3660 225564
rect 3620 201929 3648 225558
rect 3606 201920 3662 201929
rect 3606 201855 3662 201864
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3516 150408 3568 150414
rect 3516 150350 3568 150356
rect 3528 149841 3556 150350
rect 3514 149832 3570 149841
rect 3514 149767 3570 149776
rect 4816 137018 4844 257314
rect 7576 238746 7604 267106
rect 11716 244254 11744 292538
rect 11704 244248 11756 244254
rect 11704 244190 11756 244196
rect 11152 240168 11204 240174
rect 11152 240110 11204 240116
rect 7564 238740 7616 238746
rect 7564 238682 7616 238688
rect 11164 235958 11192 240110
rect 11152 235952 11204 235958
rect 11152 235894 11204 235900
rect 11704 175976 11756 175982
rect 11704 175918 11756 175924
rect 4804 137012 4856 137018
rect 4804 136954 4856 136960
rect 11716 111790 11744 175918
rect 14476 164218 14504 294578
rect 21364 289876 21416 289882
rect 21364 289818 21416 289824
rect 18604 264240 18656 264246
rect 18604 264182 18656 264188
rect 17224 229764 17276 229770
rect 17224 229706 17276 229712
rect 15844 188556 15896 188562
rect 15844 188498 15896 188504
rect 14464 164212 14516 164218
rect 14464 164154 14516 164160
rect 11704 111784 11756 111790
rect 11704 111726 11756 111732
rect 3516 97980 3568 97986
rect 3516 97922 3568 97928
rect 3528 97617 3556 97922
rect 3514 97608 3570 97617
rect 3514 97543 3570 97552
rect 3516 85536 3568 85542
rect 3516 85478 3568 85484
rect 3528 84697 3556 85478
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 4160 68332 4212 68338
rect 4160 68274 4212 68280
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 2778 36544 2834 36553
rect 2778 36479 2834 36488
rect 1308 34468 1360 34474
rect 1308 34410 1360 34416
rect 1320 33182 1348 34410
rect 20 33176 72 33182
rect 20 33118 72 33124
rect 1308 33176 1360 33182
rect 1308 33118 1360 33124
rect 32 16574 60 33118
rect 32 16546 152 16574
rect 124 354 152 16546
rect 2792 6914 2820 36479
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 2872 29708 2924 29714
rect 2872 29650 2924 29656
rect 2884 16574 2912 29650
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4172 16574 4200 68274
rect 13820 66904 13872 66910
rect 13820 66846 13872 66852
rect 12440 60036 12492 60042
rect 12440 59978 12492 59984
rect 11060 40724 11112 40730
rect 11060 40666 11112 40672
rect 6920 37936 6972 37942
rect 6920 37878 6972 37884
rect 4804 35216 4856 35222
rect 4804 35158 4856 35164
rect 2884 16546 3648 16574
rect 4172 16546 4752 16574
rect 2792 6886 2912 6914
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 1688 480 1716 3538
rect 2884 480 2912 6886
rect 542 354 654 480
rect 124 326 654 354
rect 542 -960 654 326
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3620 354 3648 16546
rect 4068 7608 4120 7614
rect 4068 7550 4120 7556
rect 4080 6497 4108 7550
rect 4066 6488 4122 6497
rect 4066 6423 4122 6432
rect 4724 3482 4752 16546
rect 4816 3602 4844 35158
rect 6932 16574 6960 37878
rect 8300 28280 8352 28286
rect 8300 28222 8352 28228
rect 8312 16574 8340 28222
rect 6932 16546 7696 16574
rect 8312 16546 8800 16574
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 4724 3454 5304 3482
rect 5276 480 5304 3454
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 6472 480 6500 3402
rect 7668 480 7696 16546
rect 8772 480 8800 16546
rect 9678 13016 9734 13025
rect 9678 12951 9734 12960
rect 4038 354 4150 480
rect 3620 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 12951
rect 11072 3534 11100 40666
rect 11152 36576 11204 36582
rect 11152 36518 11204 36524
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 11164 480 11192 36518
rect 12452 16574 12480 59978
rect 13832 16574 13860 66846
rect 15856 45558 15884 188498
rect 17236 97986 17264 229706
rect 18616 215286 18644 264182
rect 18604 215280 18656 215286
rect 18604 215222 18656 215228
rect 21376 150414 21404 289818
rect 25504 279472 25556 279478
rect 25504 279414 25556 279420
rect 21364 150408 21416 150414
rect 21364 150350 21416 150356
rect 17224 97980 17276 97986
rect 17224 97922 17276 97928
rect 22098 53136 22154 53145
rect 22098 53071 22154 53080
rect 16580 51740 16632 51746
rect 16580 51682 16632 51688
rect 15844 45552 15896 45558
rect 15844 45494 15896 45500
rect 16592 16574 16620 51682
rect 17960 49020 18012 49026
rect 17960 48962 18012 48968
rect 12452 16546 13584 16574
rect 13832 16546 14320 16574
rect 16592 16546 17080 16574
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11992 354 12020 3470
rect 13556 480 13584 16546
rect 12318 354 12430 480
rect 11992 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 15198 4856 15254 4865
rect 15198 4791 15254 4800
rect 15212 3466 15240 4791
rect 15200 3460 15252 3466
rect 15200 3402 15252 3408
rect 15936 2100 15988 2106
rect 15936 2042 15988 2048
rect 15948 480 15976 2042
rect 17052 480 17080 16546
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 48962
rect 20720 47592 20772 47598
rect 20720 47534 20772 47540
rect 19340 22772 19392 22778
rect 19340 22714 19392 22720
rect 19352 16574 19380 22714
rect 20732 16574 20760 47534
rect 22112 16574 22140 53071
rect 23480 39364 23532 39370
rect 23480 39306 23532 39312
rect 23492 16574 23520 39306
rect 19352 16546 20208 16574
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 23492 16546 24256 16574
rect 19432 6180 19484 6186
rect 19432 6122 19484 6128
rect 19444 480 19472 6122
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20180 354 20208 16546
rect 21836 480 21864 16546
rect 20598 354 20710 480
rect 20180 326 20710 354
rect 20598 -960 20710 326
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 24228 480 24256 16546
rect 25516 7614 25544 279414
rect 34348 258058 34376 379646
rect 34428 361616 34480 361622
rect 34428 361558 34480 361564
rect 34336 258052 34388 258058
rect 34336 257994 34388 258000
rect 34348 257378 34376 257994
rect 34336 257372 34388 257378
rect 34336 257314 34388 257320
rect 30380 54528 30432 54534
rect 30380 54470 30432 54476
rect 27620 50380 27672 50386
rect 27620 50322 27672 50328
rect 26240 44872 26292 44878
rect 26240 44814 26292 44820
rect 25504 7608 25556 7614
rect 25504 7550 25556 7556
rect 25320 3528 25372 3534
rect 25320 3470 25372 3476
rect 25332 480 25360 3470
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 44814
rect 27632 6914 27660 50322
rect 29000 43444 29052 43450
rect 29000 43386 29052 43392
rect 27712 42152 27764 42158
rect 27712 42094 27764 42100
rect 27724 16574 27752 42094
rect 29012 16574 29040 43386
rect 30392 16574 30420 54470
rect 31760 47660 31812 47666
rect 31760 47602 31812 47608
rect 31772 16574 31800 47602
rect 33140 42084 33192 42090
rect 33140 42026 33192 42032
rect 33152 16574 33180 42026
rect 34440 21418 34468 361558
rect 35268 336734 35296 474710
rect 40052 387122 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 57244 702500 57296 702506
rect 57244 702442 57296 702448
rect 42800 400920 42852 400926
rect 42800 400862 42852 400868
rect 42812 400246 42840 400862
rect 42800 400240 42852 400246
rect 42800 400182 42852 400188
rect 44088 400240 44140 400246
rect 44088 400182 44140 400188
rect 40868 399492 40920 399498
rect 40868 399434 40920 399440
rect 40880 398886 40908 399434
rect 40868 398880 40920 398886
rect 40868 398822 40920 398828
rect 41328 398880 41380 398886
rect 41328 398822 41380 398828
rect 40040 387116 40092 387122
rect 40040 387058 40092 387064
rect 39948 376848 40000 376854
rect 39948 376790 40000 376796
rect 35808 376780 35860 376786
rect 35808 376722 35860 376728
rect 35256 336728 35308 336734
rect 35256 336670 35308 336676
rect 34888 255264 34940 255270
rect 34888 255206 34940 255212
rect 34900 254590 34928 255206
rect 35820 254590 35848 376722
rect 39304 371272 39356 371278
rect 39304 371214 39356 371220
rect 37188 367124 37240 367130
rect 37188 367066 37240 367072
rect 37096 358828 37148 358834
rect 37096 358770 37148 358776
rect 34888 254584 34940 254590
rect 34888 254526 34940 254532
rect 35808 254584 35860 254590
rect 35808 254526 35860 254532
rect 37108 235958 37136 358770
rect 37096 235952 37148 235958
rect 37096 235894 37148 235900
rect 34520 55888 34572 55894
rect 34520 55830 34572 55836
rect 34428 21412 34480 21418
rect 34428 21354 34480 21360
rect 27724 16546 28488 16574
rect 29012 16546 30144 16574
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 33152 16546 33640 16574
rect 27632 6886 27752 6914
rect 27724 480 27752 6886
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28460 354 28488 16546
rect 30116 480 30144 16546
rect 28878 354 28990 480
rect 28460 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 33612 480 33640 16546
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 55830
rect 35900 44940 35952 44946
rect 35900 44882 35952 44888
rect 35912 6914 35940 44882
rect 37200 32434 37228 367066
rect 39316 332586 39344 371214
rect 39304 332580 39356 332586
rect 39304 332522 39356 332528
rect 39856 329180 39908 329186
rect 39856 329122 39908 329128
rect 39868 244254 39896 329122
rect 39856 244248 39908 244254
rect 39856 244190 39908 244196
rect 37280 57248 37332 57254
rect 37280 57190 37332 57196
rect 37188 32428 37240 32434
rect 37188 32370 37240 32376
rect 35992 18692 36044 18698
rect 35992 18634 36044 18640
rect 36004 16574 36032 18634
rect 37292 16574 37320 57190
rect 38660 40792 38712 40798
rect 38660 40734 38712 40740
rect 38672 16574 38700 40734
rect 36004 16546 36768 16574
rect 37292 16546 38424 16574
rect 38672 16546 39160 16574
rect 35912 6886 36032 6914
rect 36004 480 36032 6886
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 38396 480 38424 16546
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39960 7682 39988 376790
rect 40684 295656 40736 295662
rect 40684 295598 40736 295604
rect 40696 20670 40724 295598
rect 41340 267714 41368 398822
rect 43996 379568 44048 379574
rect 43996 379510 44048 379516
rect 42708 350600 42760 350606
rect 42708 350542 42760 350548
rect 42720 306338 42748 350542
rect 42708 306332 42760 306338
rect 42708 306274 42760 306280
rect 42720 305726 42748 306274
rect 42708 305720 42760 305726
rect 42708 305662 42760 305668
rect 44008 268394 44036 379510
rect 44100 274650 44128 400182
rect 48228 396772 48280 396778
rect 48228 396714 48280 396720
rect 48240 396098 48268 396714
rect 48228 396092 48280 396098
rect 48228 396034 48280 396040
rect 48136 360256 48188 360262
rect 48136 360198 48188 360204
rect 46848 353320 46900 353326
rect 46848 353262 46900 353268
rect 45468 347812 45520 347818
rect 45468 347754 45520 347760
rect 44088 274644 44140 274650
rect 44088 274586 44140 274592
rect 43996 268388 44048 268394
rect 43996 268330 44048 268336
rect 44008 268122 44036 268330
rect 43444 268116 43496 268122
rect 43444 268058 43496 268064
rect 43996 268116 44048 268122
rect 43996 268058 44048 268064
rect 41328 267708 41380 267714
rect 41328 267650 41380 267656
rect 43456 33114 43484 268058
rect 45480 234598 45508 347754
rect 46860 287054 46888 353262
rect 46768 287026 46888 287054
rect 46768 280158 46796 287026
rect 46756 280152 46808 280158
rect 46756 280094 46808 280100
rect 46768 279478 46796 280094
rect 46756 279472 46808 279478
rect 46756 279414 46808 279420
rect 48044 277500 48096 277506
rect 48044 277442 48096 277448
rect 46848 277432 46900 277438
rect 46848 277374 46900 277380
rect 45468 234592 45520 234598
rect 45468 234534 45520 234540
rect 46860 220114 46888 277374
rect 46848 220108 46900 220114
rect 46848 220050 46900 220056
rect 48056 209166 48084 277442
rect 48148 264926 48176 360198
rect 48136 264920 48188 264926
rect 48136 264862 48188 264868
rect 48148 264246 48176 264862
rect 48136 264240 48188 264246
rect 48136 264182 48188 264188
rect 48240 238678 48268 396034
rect 51080 387116 51132 387122
rect 51080 387058 51132 387064
rect 51092 386578 51120 387058
rect 51080 386572 51132 386578
rect 51080 386514 51132 386520
rect 52368 386572 52420 386578
rect 52368 386514 52420 386520
rect 49608 383784 49660 383790
rect 49608 383726 49660 383732
rect 49516 263628 49568 263634
rect 49516 263570 49568 263576
rect 48228 238672 48280 238678
rect 48228 238614 48280 238620
rect 48044 209160 48096 209166
rect 48044 209102 48096 209108
rect 49528 206281 49556 263570
rect 49620 249762 49648 383726
rect 50988 381064 51040 381070
rect 50988 381006 51040 381012
rect 50896 380928 50948 380934
rect 50896 380870 50948 380876
rect 50804 276140 50856 276146
rect 50804 276082 50856 276088
rect 49608 249756 49660 249762
rect 49608 249698 49660 249704
rect 49514 206272 49570 206281
rect 49514 206207 49570 206216
rect 50816 203590 50844 276082
rect 50908 263566 50936 380870
rect 50896 263560 50948 263566
rect 50896 263502 50948 263508
rect 51000 238649 51028 381006
rect 51080 344344 51132 344350
rect 51080 344286 51132 344292
rect 51092 343670 51120 344286
rect 51080 343664 51132 343670
rect 51080 343606 51132 343612
rect 52184 343664 52236 343670
rect 52184 343606 52236 343612
rect 52196 300218 52224 343606
rect 52276 331900 52328 331906
rect 52276 331842 52328 331848
rect 52184 300212 52236 300218
rect 52184 300154 52236 300160
rect 52184 280220 52236 280226
rect 52184 280162 52236 280168
rect 50986 238640 51042 238649
rect 50986 238575 51042 238584
rect 52196 211857 52224 280162
rect 52288 235754 52316 331842
rect 52380 238814 52408 386514
rect 55128 382424 55180 382430
rect 55128 382366 55180 382372
rect 53656 379636 53708 379642
rect 53656 379578 53708 379584
rect 53564 334620 53616 334626
rect 53564 334562 53616 334568
rect 53104 293344 53156 293350
rect 53104 293286 53156 293292
rect 52368 238808 52420 238814
rect 52368 238750 52420 238756
rect 52276 235748 52328 235754
rect 52276 235690 52328 235696
rect 52182 211848 52238 211857
rect 52182 211783 52238 211792
rect 50804 203584 50856 203590
rect 50804 203526 50856 203532
rect 46940 71052 46992 71058
rect 46940 70994 46992 71000
rect 44180 61396 44232 61402
rect 44180 61338 44232 61344
rect 43444 33108 43496 33114
rect 43444 33050 43496 33056
rect 43444 29640 43496 29646
rect 43444 29582 43496 29588
rect 40684 20664 40736 20670
rect 40684 20606 40736 20612
rect 40224 14544 40276 14550
rect 40224 14486 40276 14492
rect 39948 7676 40000 7682
rect 39948 7618 40000 7624
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 14486
rect 41880 8968 41932 8974
rect 41880 8910 41932 8916
rect 41892 480 41920 8910
rect 43456 3534 43484 29582
rect 44192 3534 44220 61338
rect 45560 38004 45612 38010
rect 45560 37946 45612 37952
rect 45572 16574 45600 37946
rect 46952 16574 46980 70994
rect 49698 62792 49754 62801
rect 49698 62727 49754 62736
rect 49712 16574 49740 62727
rect 53116 59362 53144 293286
rect 53576 266354 53604 334562
rect 53668 294642 53696 379578
rect 53748 374060 53800 374066
rect 53748 374002 53800 374008
rect 53656 294636 53708 294642
rect 53656 294578 53708 294584
rect 53656 269136 53708 269142
rect 53656 269078 53708 269084
rect 53564 266348 53616 266354
rect 53564 266290 53616 266296
rect 53564 260908 53616 260914
rect 53564 260850 53616 260856
rect 53576 181490 53604 260850
rect 53564 181484 53616 181490
rect 53564 181426 53616 181432
rect 53668 178673 53696 269078
rect 53760 235822 53788 374002
rect 55036 356108 55088 356114
rect 55036 356050 55088 356056
rect 54944 344344 54996 344350
rect 54944 344286 54996 344292
rect 54760 269204 54812 269210
rect 54760 269146 54812 269152
rect 54484 253904 54536 253910
rect 54484 253846 54536 253852
rect 53748 235816 53800 235822
rect 53748 235758 53800 235764
rect 53654 178664 53710 178673
rect 53654 178599 53710 178608
rect 54496 85542 54524 253846
rect 54772 195430 54800 269146
rect 54956 267646 54984 344286
rect 54944 267640 54996 267646
rect 54944 267582 54996 267588
rect 54852 260976 54904 260982
rect 54852 260918 54904 260924
rect 54864 213246 54892 260918
rect 55048 238513 55076 356050
rect 55140 255270 55168 382366
rect 56416 382356 56468 382362
rect 56416 382298 56468 382304
rect 56324 334892 56376 334898
rect 56324 334834 56376 334840
rect 56232 264988 56284 264994
rect 56232 264930 56284 264936
rect 55128 255264 55180 255270
rect 55128 255206 55180 255212
rect 55034 238504 55090 238513
rect 55034 238439 55090 238448
rect 56244 221474 56272 264930
rect 56336 254658 56364 334834
rect 56428 293350 56456 382298
rect 57256 374066 57284 702442
rect 72988 702434 73016 703520
rect 79324 703044 79376 703050
rect 79324 702986 79376 702992
rect 71976 702406 73016 702434
rect 66168 700324 66220 700330
rect 66168 700266 66220 700272
rect 58624 670744 58676 670750
rect 58624 670686 58676 670692
rect 57796 385144 57848 385150
rect 57796 385086 57848 385092
rect 57244 374060 57296 374066
rect 57244 374002 57296 374008
rect 56508 357468 56560 357474
rect 56508 357410 56560 357416
rect 56416 293344 56468 293350
rect 56416 293286 56468 293292
rect 56416 258120 56468 258126
rect 56416 258062 56468 258068
rect 56324 254652 56376 254658
rect 56324 254594 56376 254600
rect 56232 221468 56284 221474
rect 56232 221410 56284 221416
rect 56428 214674 56456 258062
rect 56520 253910 56548 357410
rect 57704 334824 57756 334830
rect 57704 334766 57756 334772
rect 56508 253904 56560 253910
rect 56508 253846 56560 253852
rect 56508 251252 56560 251258
rect 56508 251194 56560 251200
rect 56416 214668 56468 214674
rect 56416 214610 56468 214616
rect 54852 213240 54904 213246
rect 54852 213182 54904 213188
rect 54760 195424 54812 195430
rect 54760 195366 54812 195372
rect 56520 189786 56548 251194
rect 57612 249824 57664 249830
rect 57612 249766 57664 249772
rect 57624 193934 57652 249766
rect 57716 238746 57744 334766
rect 57808 282878 57836 385086
rect 57888 357536 57940 357542
rect 57888 357478 57940 357484
rect 57900 330449 57928 357478
rect 58636 339318 58664 670686
rect 60740 565888 60792 565894
rect 60740 565830 60792 565836
rect 59268 382560 59320 382566
rect 59268 382502 59320 382508
rect 59176 364404 59228 364410
rect 59176 364346 59228 364352
rect 58624 339312 58676 339318
rect 58624 339254 58676 339260
rect 57886 330440 57942 330449
rect 57886 330375 57942 330384
rect 59188 319462 59216 364346
rect 59176 319456 59228 319462
rect 59176 319398 59228 319404
rect 57888 294160 57940 294166
rect 57888 294102 57940 294108
rect 57796 282872 57848 282878
rect 57796 282814 57848 282820
rect 57796 274712 57848 274718
rect 57796 274654 57848 274660
rect 57704 238740 57756 238746
rect 57704 238682 57756 238688
rect 57612 193928 57664 193934
rect 57612 193870 57664 193876
rect 56508 189780 56560 189786
rect 56508 189722 56560 189728
rect 57808 188358 57836 274654
rect 57796 188352 57848 188358
rect 57796 188294 57848 188300
rect 54484 85536 54536 85542
rect 54484 85478 54536 85484
rect 56598 64152 56654 64161
rect 56598 64087 56654 64096
rect 53104 59356 53156 59362
rect 53104 59298 53156 59304
rect 52460 58676 52512 58682
rect 52460 58618 52512 58624
rect 51080 39432 51132 39438
rect 51080 39374 51132 39380
rect 45572 16546 46704 16574
rect 46952 16546 47440 16574
rect 49712 16546 50200 16574
rect 44272 10328 44324 10334
rect 44272 10270 44324 10276
rect 43444 3528 43496 3534
rect 43444 3470 43496 3476
rect 44180 3528 44232 3534
rect 44180 3470 44232 3476
rect 43076 3460 43128 3466
rect 43076 3402 43128 3408
rect 43088 480 43116 3402
rect 44284 480 44312 10270
rect 45100 3528 45152 3534
rect 45100 3470 45152 3476
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45112 354 45140 3470
rect 46676 480 46704 16546
rect 45438 354 45550 480
rect 45112 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 48504 15904 48556 15910
rect 48504 15846 48556 15852
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 15846
rect 50172 480 50200 16546
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51092 354 51120 39374
rect 52472 3534 52500 58618
rect 55220 18624 55272 18630
rect 55220 18566 55272 18572
rect 55232 16574 55260 18566
rect 56612 16574 56640 64087
rect 57900 35902 57928 294102
rect 59280 280090 59308 382502
rect 60648 382492 60700 382498
rect 60648 382434 60700 382440
rect 60464 368552 60516 368558
rect 60464 368494 60516 368500
rect 60476 336122 60504 368494
rect 60556 354816 60608 354822
rect 60556 354758 60608 354764
rect 60464 336116 60516 336122
rect 60464 336058 60516 336064
rect 60464 298784 60516 298790
rect 60464 298726 60516 298732
rect 59268 280084 59320 280090
rect 59268 280026 59320 280032
rect 60280 271992 60332 271998
rect 60280 271934 60332 271940
rect 59268 271924 59320 271930
rect 59268 271866 59320 271872
rect 59084 262268 59136 262274
rect 59084 262210 59136 262216
rect 58624 254584 58676 254590
rect 58624 254526 58676 254532
rect 58636 235890 58664 254526
rect 58624 235884 58676 235890
rect 58624 235826 58676 235832
rect 59096 204950 59124 262210
rect 59176 249688 59228 249694
rect 59176 249630 59228 249636
rect 59084 204944 59136 204950
rect 59084 204886 59136 204892
rect 59188 181558 59216 249630
rect 59280 191214 59308 271866
rect 60188 230444 60240 230450
rect 60188 230386 60240 230392
rect 60200 229770 60228 230386
rect 60188 229764 60240 229770
rect 60188 229706 60240 229712
rect 60292 198150 60320 271934
rect 60372 258188 60424 258194
rect 60372 258130 60424 258136
rect 60384 218657 60412 258130
rect 60476 230450 60504 298726
rect 60568 271862 60596 354758
rect 60660 284306 60688 382434
rect 60752 345030 60780 565830
rect 65984 389292 66036 389298
rect 65984 389234 66036 389240
rect 62028 383716 62080 383722
rect 62028 383658 62080 383664
rect 61844 360324 61896 360330
rect 61844 360266 61896 360272
rect 60740 345024 60792 345030
rect 60740 344966 60792 344972
rect 60752 344350 60780 344966
rect 60740 344344 60792 344350
rect 60740 344286 60792 344292
rect 61856 316810 61884 360266
rect 61936 351960 61988 351966
rect 61936 351902 61988 351908
rect 61948 334694 61976 351902
rect 61936 334688 61988 334694
rect 61936 334630 61988 334636
rect 61936 330608 61988 330614
rect 61936 330550 61988 330556
rect 61844 316804 61896 316810
rect 61844 316746 61896 316752
rect 61844 305788 61896 305794
rect 61844 305730 61896 305736
rect 60648 284300 60700 284306
rect 60648 284242 60700 284248
rect 60556 271856 60608 271862
rect 60556 271798 60608 271804
rect 61752 270564 61804 270570
rect 61752 270506 61804 270512
rect 61384 259480 61436 259486
rect 61384 259422 61436 259428
rect 60648 257372 60700 257378
rect 60648 257314 60700 257320
rect 60464 230444 60516 230450
rect 60464 230386 60516 230392
rect 60370 218648 60426 218657
rect 60370 218583 60426 218592
rect 60280 198144 60332 198150
rect 60280 198086 60332 198092
rect 59268 191208 59320 191214
rect 59268 191150 59320 191156
rect 60660 182889 60688 257314
rect 61396 249694 61424 259422
rect 61660 254652 61712 254658
rect 61660 254594 61712 254600
rect 61672 254017 61700 254594
rect 61658 254008 61714 254017
rect 61658 253943 61714 253952
rect 61384 249688 61436 249694
rect 61384 249630 61436 249636
rect 61764 239465 61792 270506
rect 61856 245614 61884 305730
rect 61948 260846 61976 330550
rect 62040 294642 62068 383658
rect 64788 375420 64840 375426
rect 64788 375362 64840 375368
rect 63408 365764 63460 365770
rect 63408 365706 63460 365712
rect 63316 364472 63368 364478
rect 63316 364414 63368 364420
rect 63132 314084 63184 314090
rect 63132 314026 63184 314032
rect 62028 294636 62080 294642
rect 62028 294578 62080 294584
rect 61936 260840 61988 260846
rect 61936 260782 61988 260788
rect 62028 247172 62080 247178
rect 62028 247114 62080 247120
rect 61936 247104 61988 247110
rect 61936 247046 61988 247052
rect 61844 245608 61896 245614
rect 61844 245550 61896 245556
rect 61750 239456 61806 239465
rect 61750 239391 61806 239400
rect 61948 210526 61976 247046
rect 61936 210520 61988 210526
rect 61936 210462 61988 210468
rect 62040 191146 62068 247114
rect 63144 238610 63172 314026
rect 63328 300150 63356 364414
rect 63420 313954 63448 365706
rect 64604 354748 64656 354754
rect 64604 354690 64656 354696
rect 64616 316878 64644 354690
rect 64696 347880 64748 347886
rect 64696 347822 64748 347828
rect 64604 316872 64656 316878
rect 64604 316814 64656 316820
rect 63408 313948 63460 313954
rect 63408 313890 63460 313896
rect 63316 300144 63368 300150
rect 63316 300086 63368 300092
rect 64708 297401 64736 347822
rect 64694 297392 64750 297401
rect 64694 297327 64750 297336
rect 64604 274780 64656 274786
rect 64604 274722 64656 274728
rect 63316 257440 63368 257446
rect 63316 257382 63368 257388
rect 63224 256760 63276 256766
rect 63224 256702 63276 256708
rect 63236 239426 63264 256702
rect 63224 239420 63276 239426
rect 63224 239362 63276 239368
rect 63132 238604 63184 238610
rect 63132 238546 63184 238552
rect 62028 191140 62080 191146
rect 62028 191082 62080 191088
rect 63328 182986 63356 257382
rect 64512 252612 64564 252618
rect 64512 252554 64564 252560
rect 63408 241528 63460 241534
rect 63408 241470 63460 241476
rect 63420 227050 63448 241470
rect 64524 239494 64552 252554
rect 64512 239488 64564 239494
rect 64512 239430 64564 239436
rect 64616 231198 64644 274722
rect 64696 251320 64748 251326
rect 64696 251262 64748 251268
rect 64604 231192 64656 231198
rect 64604 231134 64656 231140
rect 63408 227044 63460 227050
rect 63408 226986 63460 226992
rect 64708 184210 64736 251262
rect 64696 184204 64748 184210
rect 64696 184146 64748 184152
rect 63316 182980 63368 182986
rect 63316 182922 63368 182928
rect 60646 182880 60702 182889
rect 60646 182815 60702 182824
rect 59176 181552 59228 181558
rect 59176 181494 59228 181500
rect 59268 125656 59320 125662
rect 59268 125598 59320 125604
rect 59280 95062 59308 125598
rect 62028 124228 62080 124234
rect 62028 124170 62080 124176
rect 61936 122868 61988 122874
rect 61936 122810 61988 122816
rect 59268 95056 59320 95062
rect 59268 94998 59320 95004
rect 61948 93537 61976 122810
rect 61934 93528 61990 93537
rect 61934 93463 61990 93472
rect 62040 90982 62068 124170
rect 62028 90976 62080 90982
rect 62028 90918 62080 90924
rect 60740 65544 60792 65550
rect 60740 65486 60792 65492
rect 57888 35896 57940 35902
rect 57888 35838 57940 35844
rect 57900 35222 57928 35838
rect 57888 35216 57940 35222
rect 57888 35158 57940 35164
rect 59360 26920 59412 26926
rect 59360 26862 59412 26868
rect 57980 25560 58032 25566
rect 57980 25502 58032 25508
rect 57992 16574 58020 25502
rect 55232 16546 56088 16574
rect 56612 16546 56824 16574
rect 57992 16546 58480 16574
rect 54944 14476 54996 14482
rect 54944 14418 54996 14424
rect 52552 10396 52604 10402
rect 52552 10338 52604 10344
rect 52460 3528 52512 3534
rect 52460 3470 52512 3476
rect 52564 480 52592 10338
rect 53380 3528 53432 3534
rect 53380 3470 53432 3476
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53392 354 53420 3470
rect 54956 480 54984 14418
rect 56060 480 56088 16546
rect 53718 354 53830 480
rect 53392 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58452 480 58480 16546
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 26862
rect 60752 16574 60780 65486
rect 63500 33788 63552 33794
rect 63500 33730 63552 33736
rect 62120 21480 62172 21486
rect 62120 21422 62172 21428
rect 62132 16574 62160 21422
rect 63512 16574 63540 33730
rect 64800 17406 64828 375362
rect 65996 372570 66024 389234
rect 66076 380112 66128 380118
rect 66076 380054 66128 380060
rect 65984 372564 66036 372570
rect 65984 372506 66036 372512
rect 65984 353388 66036 353394
rect 65984 353330 66036 353336
rect 65892 340944 65944 340950
rect 65892 340886 65944 340892
rect 65904 328438 65932 340886
rect 65996 339386 66024 353330
rect 65984 339380 66036 339386
rect 65984 339322 66036 339328
rect 66088 338026 66116 380054
rect 66180 354822 66208 700266
rect 68284 694816 68336 694822
rect 68284 694758 68336 694764
rect 67730 377088 67786 377097
rect 67730 377023 67786 377032
rect 67638 376952 67694 376961
rect 67638 376887 67694 376896
rect 67652 376854 67680 376887
rect 67640 376848 67692 376854
rect 67640 376790 67692 376796
rect 67744 376786 67772 377023
rect 67732 376780 67784 376786
rect 67732 376722 67784 376728
rect 67638 375728 67694 375737
rect 67638 375663 67694 375672
rect 67546 375592 67602 375601
rect 67546 375527 67602 375536
rect 67560 374678 67588 375527
rect 67652 375426 67680 375663
rect 67640 375420 67692 375426
rect 67640 375362 67692 375368
rect 67548 374672 67600 374678
rect 67548 374614 67600 374620
rect 67454 374368 67510 374377
rect 67454 374303 67510 374312
rect 67362 374232 67418 374241
rect 67362 374167 67418 374176
rect 67272 371272 67324 371278
rect 67272 371214 67324 371220
rect 66168 354816 66220 354822
rect 66168 354758 66220 354764
rect 66166 351928 66222 351937
rect 66166 351863 66222 351872
rect 66076 338020 66128 338026
rect 66076 337962 66128 337968
rect 65892 328432 65944 328438
rect 65892 328374 65944 328380
rect 66076 301504 66128 301510
rect 66076 301446 66128 301452
rect 65984 295452 66036 295458
rect 65984 295394 66036 295400
rect 65996 287026 66024 295394
rect 65984 287020 66036 287026
rect 65984 286962 66036 286968
rect 66088 285666 66116 301446
rect 66180 294778 66208 351863
rect 66168 294772 66220 294778
rect 66168 294714 66220 294720
rect 67284 288017 67312 371214
rect 67376 333266 67404 374167
rect 67364 333260 67416 333266
rect 67364 333202 67416 333208
rect 67468 329254 67496 374303
rect 67640 373992 67692 373998
rect 67640 373934 67692 373940
rect 67652 373833 67680 373934
rect 67638 373824 67694 373833
rect 67638 373759 67694 373768
rect 67640 372564 67692 372570
rect 67640 372506 67692 372512
rect 67652 371793 67680 372506
rect 67638 371784 67694 371793
rect 67638 371719 67694 371728
rect 67638 368928 67694 368937
rect 67638 368863 67694 368872
rect 67652 368558 67680 368863
rect 67640 368552 67692 368558
rect 67640 368494 67692 368500
rect 67638 367568 67694 367577
rect 67638 367503 67694 367512
rect 67652 367130 67680 367503
rect 67640 367124 67692 367130
rect 67640 367066 67692 367072
rect 67638 365800 67694 365809
rect 67638 365735 67640 365744
rect 67692 365735 67694 365744
rect 67640 365706 67692 365712
rect 67730 364848 67786 364857
rect 67730 364783 67786 364792
rect 67640 364472 67692 364478
rect 67638 364440 67640 364449
rect 67692 364440 67694 364449
rect 67744 364410 67772 364783
rect 67638 364375 67694 364384
rect 67732 364404 67784 364410
rect 67732 364346 67784 364352
rect 67638 362128 67694 362137
rect 67638 362063 67694 362072
rect 67652 361622 67680 362063
rect 67640 361616 67692 361622
rect 67640 361558 67692 361564
rect 67638 360360 67694 360369
rect 68296 360330 68324 694758
rect 70308 576904 70360 576910
rect 70308 576846 70360 576852
rect 68836 403640 68888 403646
rect 68836 403582 68888 403588
rect 68744 398132 68796 398138
rect 68744 398074 68796 398080
rect 68376 384192 68428 384198
rect 68376 384134 68428 384140
rect 67638 360295 67694 360304
rect 67732 360324 67784 360330
rect 67652 360262 67680 360295
rect 67732 360266 67784 360272
rect 68284 360324 68336 360330
rect 68284 360266 68336 360272
rect 67640 360256 67692 360262
rect 67640 360198 67692 360204
rect 67638 359408 67694 359417
rect 67638 359343 67694 359352
rect 67652 358834 67680 359343
rect 67744 359281 67772 360266
rect 67730 359272 67786 359281
rect 67730 359207 67786 359216
rect 67640 358828 67692 358834
rect 67640 358770 67692 358776
rect 67730 358048 67786 358057
rect 67730 357983 67786 357992
rect 67744 357542 67772 357983
rect 67732 357536 67784 357542
rect 67638 357504 67694 357513
rect 67732 357478 67784 357484
rect 67638 357439 67640 357448
rect 67692 357439 67694 357448
rect 67640 357410 67692 357416
rect 67638 356552 67694 356561
rect 67638 356487 67694 356496
rect 67652 356114 67680 356487
rect 67640 356108 67692 356114
rect 67640 356050 67692 356056
rect 67638 355328 67694 355337
rect 67638 355263 67694 355272
rect 67652 354754 67680 355263
rect 67730 354920 67786 354929
rect 67730 354855 67786 354864
rect 67744 354822 67772 354855
rect 67732 354816 67784 354822
rect 67732 354758 67784 354764
rect 67640 354748 67692 354754
rect 67640 354690 67692 354696
rect 67638 353968 67694 353977
rect 67638 353903 67694 353912
rect 67652 353326 67680 353903
rect 68098 353424 68154 353433
rect 68098 353359 68100 353368
rect 68152 353359 68154 353368
rect 68100 353330 68152 353336
rect 67640 353320 67692 353326
rect 67640 353262 67692 353268
rect 67638 352608 67694 352617
rect 67638 352543 67694 352552
rect 67652 351966 67680 352543
rect 67640 351960 67692 351966
rect 68388 351937 68416 384134
rect 68756 373994 68784 398074
rect 68848 386510 68876 403582
rect 68836 386504 68888 386510
rect 68836 386446 68888 386452
rect 68664 373966 68784 373994
rect 68664 371929 68692 373966
rect 68650 371920 68706 371929
rect 68650 371855 68706 371864
rect 68664 371278 68692 371855
rect 68652 371272 68704 371278
rect 68652 371214 68704 371220
rect 68558 363760 68614 363769
rect 68558 363695 68614 363704
rect 67640 351902 67692 351908
rect 68374 351928 68430 351937
rect 68374 351863 68430 351872
rect 67638 351112 67694 351121
rect 67638 351047 67694 351056
rect 67652 350606 67680 351047
rect 67640 350600 67692 350606
rect 67640 350542 67692 350548
rect 67730 348528 67786 348537
rect 67730 348463 67786 348472
rect 67638 348120 67694 348129
rect 67638 348055 67694 348064
rect 67652 347886 67680 348055
rect 67640 347880 67692 347886
rect 67640 347822 67692 347828
rect 67744 347818 67772 348463
rect 67732 347812 67784 347818
rect 67732 347754 67784 347760
rect 67640 345024 67692 345030
rect 67640 344966 67692 344972
rect 67652 344593 67680 344966
rect 67730 344720 67786 344729
rect 67730 344655 67786 344664
rect 67638 344584 67694 344593
rect 67638 344519 67694 344528
rect 67744 343670 67772 344655
rect 67732 343664 67784 343670
rect 67732 343606 67784 343612
rect 67638 341728 67694 341737
rect 67638 341663 67694 341672
rect 67652 340950 67680 341663
rect 67640 340944 67692 340950
rect 67640 340886 67692 340892
rect 68572 338774 68600 363695
rect 68848 363633 68876 386446
rect 70216 385076 70268 385082
rect 70216 385018 70268 385024
rect 70228 382566 70256 385018
rect 70216 382560 70268 382566
rect 70216 382502 70268 382508
rect 70228 379930 70256 382502
rect 70058 379902 70256 379930
rect 69110 369880 69166 369889
rect 69110 369815 69166 369824
rect 69018 368520 69074 368529
rect 69018 368455 69074 368464
rect 68834 363624 68890 363633
rect 68834 363559 68890 363568
rect 68834 349208 68890 349217
rect 68834 349143 68890 349152
rect 68742 342408 68798 342417
rect 68742 342343 68798 342352
rect 68560 338768 68612 338774
rect 68560 338710 68612 338716
rect 68756 334626 68784 342343
rect 68848 336190 68876 349143
rect 68926 340232 68982 340241
rect 68926 340167 68982 340176
rect 68836 336184 68888 336190
rect 68836 336126 68888 336132
rect 68744 334620 68796 334626
rect 68744 334562 68796 334568
rect 67456 329248 67508 329254
rect 67456 329190 67508 329196
rect 68940 322250 68968 340167
rect 68928 322244 68980 322250
rect 68928 322186 68980 322192
rect 69032 308514 69060 368455
rect 69124 329118 69152 369815
rect 69202 349888 69258 349897
rect 69202 349823 69258 349832
rect 69112 329112 69164 329118
rect 69112 329054 69164 329060
rect 69216 325145 69244 349823
rect 70320 345953 70348 576846
rect 71044 395344 71096 395350
rect 71044 395286 71096 395292
rect 70400 389224 70452 389230
rect 70400 389166 70452 389172
rect 70412 379930 70440 389166
rect 71056 383790 71084 395286
rect 71044 383784 71096 383790
rect 71044 383726 71096 383732
rect 71056 379930 71084 383726
rect 71976 380118 72004 702406
rect 75184 683188 75236 683194
rect 75184 683130 75236 683136
rect 72424 418192 72476 418198
rect 72424 418134 72476 418140
rect 72436 384198 72464 418134
rect 75000 390584 75052 390590
rect 75000 390526 75052 390532
rect 73712 386436 73764 386442
rect 73712 386378 73764 386384
rect 72424 384192 72476 384198
rect 72424 384134 72476 384140
rect 73068 383852 73120 383858
rect 73068 383794 73120 383800
rect 72974 382392 73030 382401
rect 72974 382327 73030 382336
rect 72056 382288 72108 382294
rect 72056 382230 72108 382236
rect 71964 380112 72016 380118
rect 71964 380054 72016 380060
rect 72068 379930 72096 382230
rect 72988 379930 73016 382327
rect 73080 382294 73108 383794
rect 73068 382288 73120 382294
rect 73068 382230 73120 382236
rect 70412 379902 70702 379930
rect 71056 379902 71346 379930
rect 71990 379902 72096 379930
rect 72634 379902 73016 379930
rect 71688 379772 71740 379778
rect 71688 379714 71740 379720
rect 71700 379681 71728 379714
rect 71686 379672 71742 379681
rect 71686 379607 71742 379616
rect 73724 379438 73752 386378
rect 74816 382424 74868 382430
rect 74816 382366 74868 382372
rect 74262 381168 74318 381177
rect 74262 381103 74318 381112
rect 74276 379930 74304 381103
rect 74828 379930 74856 382366
rect 74908 382220 74960 382226
rect 74908 382162 74960 382168
rect 74920 381002 74948 382162
rect 74908 380996 74960 381002
rect 74908 380938 74960 380944
rect 73922 379902 74304 379930
rect 74566 379902 74856 379930
rect 74920 379930 74948 380938
rect 75012 380066 75040 390526
rect 75196 382226 75224 683130
rect 76564 510672 76616 510678
rect 76564 510614 76616 510620
rect 76576 385082 76604 510614
rect 76656 387116 76708 387122
rect 76656 387058 76708 387064
rect 76564 385076 76616 385082
rect 76564 385018 76616 385024
rect 76668 382566 76696 387058
rect 76748 386572 76800 386578
rect 76748 386514 76800 386520
rect 76656 382560 76708 382566
rect 76656 382502 76708 382508
rect 75184 382220 75236 382226
rect 75184 382162 75236 382168
rect 75012 380038 75408 380066
rect 75380 379930 75408 380038
rect 76668 379930 76696 382502
rect 74920 379902 75210 379930
rect 75380 379902 75854 379930
rect 76498 379902 76696 379930
rect 76760 379930 76788 386514
rect 77852 382628 77904 382634
rect 77852 382570 77904 382576
rect 77864 382498 77892 382570
rect 77852 382492 77904 382498
rect 77852 382434 77904 382440
rect 77864 379930 77892 382434
rect 79336 381070 79364 702986
rect 79416 702840 79468 702846
rect 79416 702782 79468 702788
rect 79428 382634 79456 702782
rect 81348 702568 81400 702574
rect 81348 702510 81400 702516
rect 81360 385218 81388 702510
rect 89180 702434 89208 703520
rect 98644 703112 98696 703118
rect 98644 703054 98696 703060
rect 88352 702406 89208 702434
rect 86224 700392 86276 700398
rect 86224 700334 86276 700340
rect 86236 398138 86264 700334
rect 87604 670744 87656 670750
rect 87604 670686 87656 670692
rect 86224 398132 86276 398138
rect 86224 398074 86276 398080
rect 81532 393372 81584 393378
rect 81532 393314 81584 393320
rect 81348 385212 81400 385218
rect 81348 385154 81400 385160
rect 79416 382628 79468 382634
rect 79416 382570 79468 382576
rect 80704 382492 80756 382498
rect 80704 382434 80756 382440
rect 79324 381064 79376 381070
rect 79324 381006 79376 381012
rect 76760 379902 77142 379930
rect 77786 379902 77892 379930
rect 79336 379930 79364 381006
rect 80716 379930 80744 382434
rect 81360 379930 81388 385154
rect 81544 383654 81572 393314
rect 85672 387864 85724 387870
rect 85672 387806 85724 387812
rect 84936 386368 84988 386374
rect 84936 386310 84988 386316
rect 84948 383722 84976 386310
rect 84936 383716 84988 383722
rect 84936 383658 84988 383664
rect 79336 379902 79718 379930
rect 80362 379902 80744 379930
rect 81006 379902 81388 379930
rect 81452 383626 81572 383654
rect 81452 379794 81480 383626
rect 84568 382968 84620 382974
rect 84568 382910 84620 382916
rect 81900 382356 81952 382362
rect 81900 382298 81952 382304
rect 81912 379930 81940 382298
rect 83278 381304 83334 381313
rect 83278 381239 83334 381248
rect 83292 379930 83320 381239
rect 84580 379930 84608 382910
rect 84948 379930 84976 383658
rect 85304 382356 85356 382362
rect 85304 382298 85356 382304
rect 81912 379902 82294 379930
rect 82938 379902 83320 379930
rect 84226 379902 84608 379930
rect 84870 379902 84976 379930
rect 85316 379794 85344 382298
rect 85684 379930 85712 387806
rect 87616 386374 87644 670686
rect 88352 388482 88380 702406
rect 93124 501016 93176 501022
rect 93124 500958 93176 500964
rect 90364 453348 90416 453354
rect 90364 453290 90416 453296
rect 89720 398880 89772 398886
rect 89720 398822 89772 398828
rect 88340 388476 88392 388482
rect 88340 388418 88392 388424
rect 87604 386368 87656 386374
rect 87604 386310 87656 386316
rect 88248 385348 88300 385354
rect 88248 385290 88300 385296
rect 87696 382560 87748 382566
rect 87696 382502 87748 382508
rect 87708 379930 87736 382502
rect 88260 379930 88288 385290
rect 89626 383752 89682 383761
rect 89626 383687 89682 383696
rect 89640 379930 89668 383687
rect 85684 379902 86158 379930
rect 87446 379902 87736 379930
rect 88090 379902 88288 379930
rect 89378 379902 89668 379930
rect 89732 379930 89760 398822
rect 90376 385286 90404 453290
rect 91744 399492 91796 399498
rect 91744 399434 91796 399440
rect 90364 385280 90416 385286
rect 90364 385222 90416 385228
rect 89812 382424 89864 382430
rect 89812 382366 89864 382372
rect 89824 380225 89852 382366
rect 89810 380216 89866 380225
rect 89810 380151 89866 380160
rect 90376 379930 90404 385222
rect 91756 383897 91784 399434
rect 93136 383926 93164 500958
rect 97264 456816 97316 456822
rect 97264 456758 97316 456764
rect 97276 399498 97304 456758
rect 97356 404388 97408 404394
rect 97356 404330 97408 404336
rect 97264 399492 97316 399498
rect 97264 399434 97316 399440
rect 94686 387832 94742 387841
rect 94686 387767 94742 387776
rect 94596 385076 94648 385082
rect 94596 385018 94648 385024
rect 93124 383920 93176 383926
rect 91742 383888 91798 383897
rect 93124 383862 93176 383868
rect 91742 383823 91798 383832
rect 91558 381032 91614 381041
rect 91558 380967 91614 380976
rect 91572 379930 91600 380967
rect 89732 379902 90022 379930
rect 90376 379902 90666 379930
rect 91310 379902 91600 379930
rect 91756 379930 91784 383823
rect 93136 383654 93164 383862
rect 93044 383626 93164 383654
rect 92848 382424 92900 382430
rect 92848 382366 92900 382372
rect 92860 379930 92888 382366
rect 91756 379902 91954 379930
rect 92598 379902 92888 379930
rect 93044 379794 93072 383626
rect 94608 379930 94636 385018
rect 94530 379902 94636 379930
rect 94700 379930 94728 387767
rect 97368 387122 97396 404330
rect 97356 387116 97408 387122
rect 97356 387058 97408 387064
rect 98656 385150 98684 703054
rect 101404 514820 101456 514826
rect 101404 514762 101456 514768
rect 99380 400240 99432 400246
rect 99380 400182 99432 400188
rect 98644 385144 98696 385150
rect 98644 385086 98696 385092
rect 96528 383988 96580 383994
rect 96528 383930 96580 383936
rect 96160 382628 96212 382634
rect 96160 382570 96212 382576
rect 96172 379930 96200 382570
rect 96540 379930 96568 383930
rect 97908 383784 97960 383790
rect 97908 383726 97960 383732
rect 97448 381132 97500 381138
rect 97448 381074 97500 381080
rect 97460 379930 97488 381074
rect 97920 379930 97948 383726
rect 98656 379930 98684 385086
rect 94700 379902 95174 379930
rect 95818 379902 96200 379930
rect 96462 379902 96568 379930
rect 97106 379902 97488 379930
rect 97750 379902 97948 379930
rect 98394 379902 98684 379930
rect 99392 379930 99420 400182
rect 101416 386578 101444 514762
rect 102140 387932 102192 387938
rect 102140 387874 102192 387880
rect 100760 386572 100812 386578
rect 100760 386514 100812 386520
rect 101404 386572 101456 386578
rect 101404 386514 101456 386520
rect 100668 385144 100720 385150
rect 100668 385086 100720 385092
rect 100680 382974 100708 385086
rect 100668 382968 100720 382974
rect 100668 382910 100720 382916
rect 100772 379930 100800 386514
rect 102152 383654 102180 387874
rect 104912 387802 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 106280 702976 106332 702982
rect 106280 702918 106332 702924
rect 104900 387796 104952 387802
rect 104900 387738 104952 387744
rect 103888 383716 103940 383722
rect 103888 383658 103940 383664
rect 102152 383626 102364 383654
rect 101864 382696 101916 382702
rect 101864 382638 101916 382644
rect 101876 379930 101904 382638
rect 102336 379930 102364 383626
rect 103900 379930 103928 383658
rect 104808 382356 104860 382362
rect 104808 382298 104860 382304
rect 104624 381064 104676 381070
rect 104624 381006 104676 381012
rect 99392 379902 99682 379930
rect 100772 379902 100970 379930
rect 101614 379902 101904 379930
rect 102258 379902 102364 379930
rect 103546 379902 103928 379930
rect 104636 379794 104664 381006
rect 104820 380186 104848 382298
rect 106188 382288 106240 382294
rect 106188 382230 106240 382236
rect 104808 380180 104860 380186
rect 104808 380122 104860 380128
rect 106200 379930 106228 382230
rect 106122 379902 106228 379930
rect 81452 379766 81650 379794
rect 85316 379766 85514 379794
rect 93044 379766 93242 379794
rect 104636 379766 104834 379794
rect 78772 379704 78824 379710
rect 78824 379652 79074 379658
rect 78772 379646 79074 379652
rect 78784 379630 79074 379646
rect 99944 379642 100326 379658
rect 99932 379636 100326 379642
rect 99984 379630 100326 379636
rect 102902 379642 103192 379658
rect 102902 379636 103204 379642
rect 102902 379630 103152 379636
rect 99932 379578 99984 379584
rect 103152 379578 103204 379584
rect 105084 379568 105136 379574
rect 86958 379536 87014 379545
rect 86802 379494 86958 379522
rect 106292 379522 106320 702918
rect 117228 702908 117280 702914
rect 117228 702850 117280 702856
rect 115848 702636 115900 702642
rect 115848 702578 115900 702584
rect 110420 698964 110472 698970
rect 110420 698906 110472 698912
rect 108304 422340 108356 422346
rect 108304 422282 108356 422288
rect 108316 389366 108344 422282
rect 108304 389360 108356 389366
rect 108304 389302 108356 389308
rect 109684 389360 109736 389366
rect 109684 389302 109736 389308
rect 109696 385422 109724 389302
rect 109684 385416 109736 385422
rect 109684 385358 109736 385364
rect 106832 382492 106884 382498
rect 106832 382434 106884 382440
rect 106844 380254 106872 382434
rect 106832 380248 106884 380254
rect 106832 380190 106884 380196
rect 109696 379930 109724 385358
rect 109868 382560 109920 382566
rect 109868 382502 109920 382508
rect 109776 381132 109828 381138
rect 109776 381074 109828 381080
rect 109342 379902 109724 379930
rect 109500 379772 109552 379778
rect 109500 379714 109552 379720
rect 107016 379568 107068 379574
rect 105136 379516 105478 379522
rect 105084 379510 105478 379516
rect 105096 379494 105478 379510
rect 106292 379516 107016 379522
rect 106292 379510 107068 379516
rect 106292 379494 107056 379510
rect 107410 379506 107700 379522
rect 107410 379500 107712 379506
rect 107410 379494 107660 379500
rect 86958 379471 87014 379480
rect 107660 379442 107712 379448
rect 71688 379432 71740 379438
rect 71686 379400 71688 379409
rect 73712 379432 73764 379438
rect 71740 379400 71742 379409
rect 108946 379400 109002 379409
rect 73712 379374 73764 379380
rect 108054 379358 108344 379386
rect 108698 379358 108946 379386
rect 71686 379335 71742 379344
rect 108316 379302 108344 379358
rect 108946 379335 109002 379344
rect 108304 379296 108356 379302
rect 108304 379238 108356 379244
rect 109512 379137 109540 379714
rect 109684 379500 109736 379506
rect 109684 379442 109736 379448
rect 109498 379128 109554 379137
rect 109498 379063 109554 379072
rect 109696 370530 109724 379442
rect 109788 373697 109816 381074
rect 109880 377777 109908 382502
rect 109866 377768 109922 377777
rect 109866 377703 109922 377712
rect 109774 373688 109830 373697
rect 109774 373623 109830 373632
rect 109684 370524 109736 370530
rect 109684 370466 109736 370472
rect 110326 366616 110382 366625
rect 110326 366551 110382 366560
rect 110340 365770 110368 366551
rect 109316 365764 109368 365770
rect 109316 365706 109368 365712
rect 110328 365764 110380 365770
rect 110328 365706 110380 365712
rect 109328 354674 109356 365706
rect 109592 361548 109644 361554
rect 109592 361490 109644 361496
rect 109604 360777 109632 361490
rect 109590 360768 109646 360777
rect 109590 360703 109646 360712
rect 109498 358184 109554 358193
rect 109498 358119 109554 358128
rect 109144 354646 109356 354674
rect 69294 345944 69350 345953
rect 69294 345879 69350 345888
rect 70306 345944 70362 345953
rect 70306 345879 70362 345888
rect 69308 331945 69336 345879
rect 70490 341048 70546 341057
rect 70490 340983 70546 340992
rect 70044 337006 70072 340068
rect 70504 339998 70532 340983
rect 70492 339992 70544 339998
rect 70492 339934 70544 339940
rect 70688 337754 70716 340068
rect 70676 337748 70728 337754
rect 70676 337690 70728 337696
rect 71332 337618 71360 340068
rect 71320 337612 71372 337618
rect 71320 337554 71372 337560
rect 70032 337000 70084 337006
rect 70032 336942 70084 336948
rect 69294 331936 69350 331945
rect 69294 331871 69350 331880
rect 69202 325136 69258 325145
rect 69202 325071 69258 325080
rect 71044 322380 71096 322386
rect 71044 322322 71096 322328
rect 69020 308508 69072 308514
rect 69020 308450 69072 308456
rect 67456 303680 67508 303686
rect 67456 303622 67508 303628
rect 67270 288008 67326 288017
rect 67270 287943 67326 287952
rect 67468 287881 67496 303622
rect 69020 303000 69072 303006
rect 69020 302942 69072 302948
rect 67548 296880 67600 296886
rect 67548 296822 67600 296828
rect 67560 290873 67588 296822
rect 68742 293992 68798 294001
rect 68742 293927 68798 293936
rect 68652 292596 68704 292602
rect 68652 292538 68704 292544
rect 68006 291136 68062 291145
rect 68006 291071 68062 291080
rect 67546 290864 67602 290873
rect 67546 290799 67602 290808
rect 68020 289882 68048 291071
rect 68008 289876 68060 289882
rect 68008 289818 68060 289824
rect 67546 288552 67602 288561
rect 67546 288487 67602 288496
rect 67454 287872 67510 287881
rect 67454 287807 67510 287816
rect 66076 285660 66128 285666
rect 66076 285602 66128 285608
rect 67454 276312 67510 276321
rect 67454 276247 67510 276256
rect 66168 268252 66220 268258
rect 66168 268194 66220 268200
rect 65892 249892 65944 249898
rect 65892 249834 65944 249840
rect 65904 239970 65932 249834
rect 66076 248668 66128 248674
rect 66076 248610 66128 248616
rect 65984 244316 66036 244322
rect 65984 244258 66036 244264
rect 65892 239964 65944 239970
rect 65892 239906 65944 239912
rect 65996 185910 66024 244258
rect 65984 185904 66036 185910
rect 65984 185846 66036 185852
rect 66088 180198 66116 248610
rect 66076 180192 66128 180198
rect 66076 180134 66128 180140
rect 66180 178770 66208 268194
rect 67468 185638 67496 276247
rect 67456 185632 67508 185638
rect 67456 185574 67508 185580
rect 67560 184346 67588 288487
rect 67730 287056 67786 287065
rect 67730 286991 67732 287000
rect 67784 286991 67786 287000
rect 67732 286962 67784 286968
rect 68192 285660 68244 285666
rect 68192 285602 68244 285608
rect 68204 285433 68232 285602
rect 68190 285424 68246 285433
rect 68190 285359 68246 285368
rect 68664 284753 68692 292538
rect 68756 286113 68784 293927
rect 69032 291145 69060 302942
rect 70674 296848 70730 296857
rect 70674 296783 70730 296792
rect 70032 294432 70084 294438
rect 70032 294374 70084 294380
rect 70044 291924 70072 294374
rect 70688 291963 70716 296783
rect 71056 292369 71084 322322
rect 71976 312662 72004 340068
rect 72424 337748 72476 337754
rect 72424 337690 72476 337696
rect 72436 313993 72464 337690
rect 72620 336802 72648 340068
rect 73264 337482 73292 340068
rect 73908 338026 73936 340068
rect 73896 338020 73948 338026
rect 73896 337962 73948 337968
rect 73804 337612 73856 337618
rect 73804 337554 73856 337560
rect 73252 337476 73304 337482
rect 73252 337418 73304 337424
rect 72608 336796 72660 336802
rect 72608 336738 72660 336744
rect 73160 327820 73212 327826
rect 73160 327762 73212 327768
rect 72422 313984 72478 313993
rect 72422 313919 72478 313928
rect 71964 312656 72016 312662
rect 71964 312598 72016 312604
rect 72424 311228 72476 311234
rect 72424 311170 72476 311176
rect 72240 304292 72292 304298
rect 72240 304234 72292 304240
rect 71962 298344 72018 298353
rect 71962 298279 72018 298288
rect 71320 295996 71372 296002
rect 71320 295938 71372 295944
rect 71042 292360 71098 292369
rect 71042 292295 71098 292304
rect 71332 291963 71360 295938
rect 71976 291963 72004 298279
rect 72252 291977 72280 304234
rect 72436 296002 72464 311170
rect 72424 295996 72476 296002
rect 72424 295938 72476 295944
rect 73172 294370 73200 327762
rect 73816 309777 73844 337554
rect 73908 324970 73936 337962
rect 74552 337414 74580 340068
rect 74540 337408 74592 337414
rect 74540 337350 74592 337356
rect 75276 337000 75328 337006
rect 75276 336942 75328 336948
rect 75184 336796 75236 336802
rect 75184 336738 75236 336744
rect 73896 324964 73948 324970
rect 73896 324906 73948 324912
rect 73802 309768 73858 309777
rect 73802 309703 73858 309712
rect 74540 302388 74592 302394
rect 74540 302330 74592 302336
rect 73252 300960 73304 300966
rect 73252 300902 73304 300908
rect 73160 294364 73212 294370
rect 73160 294306 73212 294312
rect 72252 291949 72634 291977
rect 73264 291963 73292 300902
rect 73620 294364 73672 294370
rect 73620 294306 73672 294312
rect 73632 291977 73660 294306
rect 73632 291949 73922 291977
rect 74552 291963 74580 302330
rect 75196 301481 75224 336738
rect 75288 309806 75316 336942
rect 75840 309874 75868 340068
rect 76484 316742 76512 340068
rect 76562 339960 76618 339969
rect 76562 339895 76618 339904
rect 76472 316736 76524 316742
rect 76472 316678 76524 316684
rect 75920 310548 75972 310554
rect 75920 310490 75972 310496
rect 75828 309868 75880 309874
rect 75828 309810 75880 309816
rect 75276 309800 75328 309806
rect 75276 309742 75328 309748
rect 75182 301472 75238 301481
rect 75182 301407 75238 301416
rect 75182 295488 75238 295497
rect 75182 295423 75238 295432
rect 75196 291963 75224 295423
rect 75826 294128 75882 294137
rect 75826 294063 75882 294072
rect 75840 291963 75868 294063
rect 75932 291977 75960 310490
rect 76576 307154 76604 339895
rect 77128 318102 77156 340068
rect 77772 337385 77800 340068
rect 78416 338026 78444 340068
rect 78404 338020 78456 338026
rect 78404 337962 78456 337968
rect 77390 337376 77446 337385
rect 77390 337311 77446 337320
rect 77758 337376 77814 337385
rect 77758 337311 77814 337320
rect 77116 318096 77168 318102
rect 77116 318038 77168 318044
rect 76564 307148 76616 307154
rect 76564 307090 76616 307096
rect 77114 293176 77170 293185
rect 77114 293111 77170 293120
rect 75932 291949 76498 291977
rect 77128 291963 77156 293111
rect 77404 291977 77432 337311
rect 79060 327758 79088 340068
rect 79324 339992 79376 339998
rect 79324 339934 79376 339940
rect 79048 327752 79100 327758
rect 79048 327694 79100 327700
rect 79336 319530 79364 339934
rect 79324 319524 79376 319530
rect 79324 319466 79376 319472
rect 79704 311166 79732 340068
rect 80992 337958 81020 340068
rect 80980 337952 81032 337958
rect 80980 337894 81032 337900
rect 80428 337476 80480 337482
rect 80428 337418 80480 337424
rect 80440 331226 80468 337418
rect 80992 336025 81020 337894
rect 81636 337482 81664 340068
rect 82280 337521 82308 340068
rect 82266 337512 82322 337521
rect 81624 337476 81676 337482
rect 82266 337447 82322 337456
rect 81624 337418 81676 337424
rect 80978 336016 81034 336025
rect 80978 335951 81034 335960
rect 82924 334898 82952 340068
rect 83568 339454 83596 340068
rect 83556 339448 83608 339454
rect 83556 339390 83608 339396
rect 83568 335354 83596 339390
rect 84212 337890 84240 340068
rect 84856 339454 84884 340068
rect 84844 339448 84896 339454
rect 84844 339390 84896 339396
rect 84200 337884 84252 337890
rect 84200 337826 84252 337832
rect 83476 335326 83596 335354
rect 82912 334892 82964 334898
rect 82912 334834 82964 334840
rect 80428 331220 80480 331226
rect 80428 331162 80480 331168
rect 79692 311160 79744 311166
rect 79692 311102 79744 311108
rect 80060 308440 80112 308446
rect 80060 308382 80112 308388
rect 79324 303748 79376 303754
rect 79324 303690 79376 303696
rect 78404 294772 78456 294778
rect 78404 294714 78456 294720
rect 77404 291949 77786 291977
rect 78416 291963 78444 294714
rect 79048 294704 79100 294710
rect 79048 294646 79100 294652
rect 79060 291963 79088 294646
rect 79336 291938 79364 303690
rect 80072 291977 80100 308382
rect 81440 306468 81492 306474
rect 81440 306410 81492 306416
rect 81452 306374 81480 306410
rect 81452 306346 81940 306374
rect 80612 299668 80664 299674
rect 80612 299610 80664 299616
rect 80152 294024 80204 294030
rect 80152 293966 80204 293972
rect 80164 293282 80192 293966
rect 80152 293276 80204 293282
rect 80152 293218 80204 293224
rect 80072 291949 80362 291977
rect 80624 291938 80652 299610
rect 81622 295352 81678 295361
rect 81622 295287 81678 295296
rect 81636 291963 81664 295287
rect 81912 291938 81940 306346
rect 83476 298858 83504 335326
rect 84292 323604 84344 323610
rect 84292 323546 84344 323552
rect 83464 298852 83516 298858
rect 83464 298794 83516 298800
rect 84200 298444 84252 298450
rect 84200 298386 84252 298392
rect 82912 295724 82964 295730
rect 82912 295666 82964 295672
rect 82924 291963 82952 295666
rect 83556 295520 83608 295526
rect 83556 295462 83608 295468
rect 83568 291963 83596 295462
rect 84212 291963 84240 298386
rect 84304 291938 84332 323546
rect 84856 314090 84884 339390
rect 84844 314084 84896 314090
rect 84844 314026 84896 314032
rect 86144 305658 86172 340068
rect 86132 305652 86184 305658
rect 86132 305594 86184 305600
rect 86788 302938 86816 340068
rect 87432 337618 87460 340068
rect 87420 337612 87472 337618
rect 87420 337554 87472 337560
rect 87604 337408 87656 337414
rect 87604 337350 87656 337356
rect 87616 325009 87644 337350
rect 87602 325000 87658 325009
rect 87602 324935 87658 324944
rect 87604 308644 87656 308650
rect 87604 308586 87656 308592
rect 86776 302932 86828 302938
rect 86776 302874 86828 302880
rect 85580 300892 85632 300898
rect 85580 300834 85632 300840
rect 85488 294976 85540 294982
rect 85488 294918 85540 294924
rect 85500 291963 85528 294918
rect 85592 291938 85620 300834
rect 87420 298376 87472 298382
rect 87420 298318 87472 298324
rect 86776 298172 86828 298178
rect 86776 298114 86828 298120
rect 86788 291963 86816 298114
rect 87432 291963 87460 298318
rect 87616 294982 87644 308586
rect 88076 307086 88104 340068
rect 88720 336054 88748 340068
rect 89076 337612 89128 337618
rect 89076 337554 89128 337560
rect 88984 336116 89036 336122
rect 88984 336058 89036 336064
rect 88708 336048 88760 336054
rect 88708 335990 88760 335996
rect 88064 307080 88116 307086
rect 88064 307022 88116 307028
rect 88340 305040 88392 305046
rect 88340 304982 88392 304988
rect 87604 294976 87656 294982
rect 87604 294918 87656 294924
rect 88352 294370 88380 304982
rect 88996 302841 89024 336058
rect 89088 308582 89116 337554
rect 89364 315314 89392 340068
rect 89352 315308 89404 315314
rect 89352 315250 89404 315256
rect 89076 308576 89128 308582
rect 89076 308518 89128 308524
rect 89720 306400 89772 306406
rect 89720 306342 89772 306348
rect 90008 306374 90036 340068
rect 91100 339312 91152 339318
rect 91100 339254 91152 339260
rect 90088 337884 90140 337890
rect 90088 337826 90140 337832
rect 90100 336122 90128 337826
rect 90088 336116 90140 336122
rect 90088 336058 90140 336064
rect 90008 306346 90220 306374
rect 88982 302832 89038 302841
rect 88982 302767 89038 302776
rect 88432 299532 88484 299538
rect 88432 299474 88484 299480
rect 88340 294364 88392 294370
rect 88340 294306 88392 294312
rect 88064 294296 88116 294302
rect 88064 294238 88116 294244
rect 88076 291963 88104 294238
rect 88444 291977 88472 299474
rect 89076 294364 89128 294370
rect 89076 294306 89128 294312
rect 89088 291977 89116 294306
rect 89732 291977 89760 306342
rect 89812 299736 89864 299742
rect 89812 299678 89864 299684
rect 89824 294352 89852 299678
rect 89824 294324 90128 294352
rect 90100 291977 90128 294324
rect 90192 293321 90220 306346
rect 91112 301617 91140 339254
rect 91296 331906 91324 340068
rect 91940 339318 91968 340068
rect 91928 339312 91980 339318
rect 91928 339254 91980 339260
rect 92584 337414 92612 340068
rect 92572 337408 92624 337414
rect 92572 337350 92624 337356
rect 91284 331900 91336 331906
rect 91284 331842 91336 331848
rect 93228 304201 93256 340068
rect 93872 322318 93900 340068
rect 94516 334830 94544 340068
rect 95160 339318 95188 340068
rect 95148 339312 95200 339318
rect 95148 339254 95200 339260
rect 94504 334824 94556 334830
rect 94504 334766 94556 334772
rect 93860 322312 93912 322318
rect 93860 322254 93912 322260
rect 95160 318782 95188 339254
rect 96448 336734 96476 340068
rect 95884 336728 95936 336734
rect 95884 336670 95936 336676
rect 96436 336728 96488 336734
rect 96436 336670 96488 336676
rect 95148 318776 95200 318782
rect 95148 318718 95200 318724
rect 94504 314016 94556 314022
rect 94504 313958 94556 313964
rect 94516 306374 94544 313958
rect 94424 306346 94544 306374
rect 93214 304192 93270 304201
rect 93214 304127 93270 304136
rect 91098 301608 91154 301617
rect 91098 301543 91154 301552
rect 93950 300112 94006 300121
rect 93950 300047 94006 300056
rect 93216 295588 93268 295594
rect 93216 295530 93268 295536
rect 92756 295180 92808 295186
rect 92756 295122 92808 295128
rect 91284 294636 91336 294642
rect 91284 294578 91336 294584
rect 90178 293312 90234 293321
rect 90178 293247 90234 293256
rect 88444 291949 88734 291977
rect 89088 291949 89378 291977
rect 89732 291949 90022 291977
rect 90100 291949 90666 291977
rect 91296 291963 91324 294578
rect 91928 294092 91980 294098
rect 91928 294034 91980 294040
rect 91940 291963 91968 294034
rect 92768 294030 92796 295122
rect 92756 294024 92808 294030
rect 92756 293966 92808 293972
rect 92768 291977 92796 293966
rect 92598 291949 92796 291977
rect 93228 291963 93256 295530
rect 93964 294370 93992 300047
rect 94424 295186 94452 306346
rect 95896 305862 95924 336670
rect 97092 323678 97120 340068
rect 97736 334665 97764 340068
rect 97722 334656 97778 334665
rect 97722 334591 97778 334600
rect 98380 330546 98408 340068
rect 98978 339810 99006 340068
rect 98656 339782 99006 339810
rect 98656 338094 98684 339782
rect 98644 338088 98696 338094
rect 98644 338030 98696 338036
rect 98368 330540 98420 330546
rect 98368 330482 98420 330488
rect 97080 323672 97132 323678
rect 97080 323614 97132 323620
rect 95884 305856 95936 305862
rect 95884 305798 95936 305804
rect 98000 300212 98052 300218
rect 98000 300154 98052 300160
rect 97356 299600 97408 299606
rect 97356 299542 97408 299548
rect 94504 297492 94556 297498
rect 94504 297434 94556 297440
rect 94412 295180 94464 295186
rect 94412 295122 94464 295128
rect 93952 294364 94004 294370
rect 93952 294306 94004 294312
rect 93860 292732 93912 292738
rect 93860 292674 93912 292680
rect 93872 291963 93900 292674
rect 94516 291963 94544 297434
rect 94780 294364 94832 294370
rect 94780 294306 94832 294312
rect 94792 291938 94820 294306
rect 96436 294228 96488 294234
rect 96436 294170 96488 294176
rect 95792 294160 95844 294166
rect 95792 294102 95844 294108
rect 95804 291963 95832 294102
rect 96448 291963 96476 294170
rect 97080 293344 97132 293350
rect 97080 293286 97132 293292
rect 97092 291963 97120 293286
rect 97368 291938 97396 299542
rect 98012 291977 98040 300154
rect 98656 297430 98684 338030
rect 99668 334762 99696 340068
rect 100312 337754 100340 340068
rect 100300 337748 100352 337754
rect 100300 337690 100352 337696
rect 101404 337748 101456 337754
rect 101404 337690 101456 337696
rect 100024 337612 100076 337618
rect 100024 337554 100076 337560
rect 99656 334756 99708 334762
rect 99656 334698 99708 334704
rect 99748 334756 99800 334762
rect 99748 334698 99800 334704
rect 99760 332586 99788 334698
rect 99748 332580 99800 332586
rect 99748 332522 99800 332528
rect 98644 297424 98696 297430
rect 98644 297366 98696 297372
rect 100036 296818 100064 337554
rect 101416 320890 101444 337690
rect 101404 320884 101456 320890
rect 101404 320826 101456 320832
rect 101404 318776 101456 318782
rect 101404 318718 101456 318724
rect 100852 302456 100904 302462
rect 100852 302398 100904 302404
rect 100024 296812 100076 296818
rect 100024 296754 100076 296760
rect 99012 296744 99064 296750
rect 99012 296686 99064 296692
rect 98012 291949 98394 291977
rect 99024 291963 99052 296686
rect 100036 294370 100064 296754
rect 100024 294364 100076 294370
rect 100024 294306 100076 294312
rect 99656 292664 99708 292670
rect 99656 292606 99708 292612
rect 99668 291963 99696 292606
rect 100864 291977 100892 302398
rect 101416 295322 101444 318718
rect 101600 308718 101628 340068
rect 102244 339425 102272 340068
rect 102230 339416 102286 339425
rect 102230 339351 102286 339360
rect 102888 329186 102916 340068
rect 102876 329180 102928 329186
rect 102876 329122 102928 329128
rect 102140 323740 102192 323746
rect 102140 323682 102192 323688
rect 102152 322386 102180 323682
rect 102140 322380 102192 322386
rect 102140 322322 102192 322328
rect 103532 311234 103560 340068
rect 104176 338094 104204 340068
rect 104164 338088 104216 338094
rect 104164 338030 104216 338036
rect 104176 333305 104204 338030
rect 104162 333296 104218 333305
rect 104162 333231 104218 333240
rect 103520 311228 103572 311234
rect 103520 311170 103572 311176
rect 101588 308712 101640 308718
rect 101588 308654 101640 308660
rect 104820 305697 104848 340068
rect 105464 327729 105492 340068
rect 106280 338904 106332 338910
rect 106280 338846 106332 338852
rect 105544 338836 105596 338842
rect 105544 338778 105596 338784
rect 105450 327720 105506 327729
rect 105450 327655 105506 327664
rect 104806 305688 104862 305697
rect 104806 305623 104862 305632
rect 103612 302252 103664 302258
rect 103612 302194 103664 302200
rect 102140 301028 102192 301034
rect 102140 300970 102192 300976
rect 101404 295316 101456 295322
rect 101404 295258 101456 295264
rect 101588 294364 101640 294370
rect 101588 294306 101640 294312
rect 100864 291949 100970 291977
rect 101600 291963 101628 294306
rect 102152 291977 102180 300970
rect 102324 299804 102376 299810
rect 102324 299746 102376 299752
rect 102152 291949 102258 291977
rect 102336 291938 102364 299746
rect 103520 292120 103572 292126
rect 103520 292062 103572 292068
rect 103532 291963 103560 292062
rect 103624 291938 103652 302194
rect 105556 298790 105584 338778
rect 106186 336696 106242 336705
rect 106186 336631 106242 336640
rect 106200 306374 106228 336631
rect 105832 306346 106228 306374
rect 105832 299577 105860 306346
rect 106096 303816 106148 303822
rect 106096 303758 106148 303764
rect 105818 299568 105874 299577
rect 105818 299503 105874 299512
rect 105544 298784 105596 298790
rect 105544 298726 105596 298732
rect 104808 295316 104860 295322
rect 104808 295258 104860 295264
rect 104820 291963 104848 295258
rect 105452 294296 105504 294302
rect 105452 294238 105504 294244
rect 105464 291963 105492 294238
rect 105832 291977 105860 299503
rect 106108 294302 106136 303758
rect 106292 294370 106320 338846
rect 106752 326398 106780 340068
rect 107396 333946 107424 340068
rect 107568 339992 107620 339998
rect 107568 339934 107620 339940
rect 107580 337958 107608 339934
rect 107994 339810 108022 340068
rect 107764 339782 108022 339810
rect 107568 337952 107620 337958
rect 107568 337894 107620 337900
rect 107384 333940 107436 333946
rect 107384 333882 107436 333888
rect 107396 332654 107424 333882
rect 107764 333878 107792 339782
rect 107752 333872 107804 333878
rect 107752 333814 107804 333820
rect 106924 332648 106976 332654
rect 106924 332590 106976 332596
rect 107384 332648 107436 332654
rect 107384 332590 107436 332596
rect 106740 326392 106792 326398
rect 106740 326334 106792 326340
rect 106936 308650 106964 332590
rect 106924 308644 106976 308650
rect 106924 308586 106976 308592
rect 106372 302320 106424 302326
rect 106372 302262 106424 302268
rect 106280 294364 106332 294370
rect 106280 294306 106332 294312
rect 106096 294296 106148 294302
rect 106096 294238 106148 294244
rect 105832 291949 106122 291977
rect 106384 291938 106412 302262
rect 107764 297498 107792 333814
rect 108684 314022 108712 340068
rect 109144 327826 109172 354646
rect 109328 337550 109356 340068
rect 109316 337544 109368 337550
rect 109316 337486 109368 337492
rect 109132 327820 109184 327826
rect 109132 327762 109184 327768
rect 109512 323610 109540 358119
rect 109604 338910 109632 360703
rect 110432 358465 110460 698906
rect 111800 530596 111852 530602
rect 111800 530538 111852 530544
rect 110604 409896 110656 409902
rect 110604 409838 110656 409844
rect 110510 378176 110566 378185
rect 110510 378111 110566 378120
rect 110418 358456 110474 358465
rect 110418 358391 110474 358400
rect 110418 340776 110474 340785
rect 110418 340711 110474 340720
rect 110328 340196 110380 340202
rect 110328 340138 110380 340144
rect 109592 338904 109644 338910
rect 109592 338846 109644 338852
rect 109500 323604 109552 323610
rect 109500 323546 109552 323552
rect 108672 314016 108724 314022
rect 108672 313958 108724 313964
rect 107752 297492 107804 297498
rect 107752 297434 107804 297440
rect 108672 296812 108724 296818
rect 108672 296754 108724 296760
rect 107108 294364 107160 294370
rect 107108 294306 107160 294312
rect 107120 291977 107148 294306
rect 107120 291949 107410 291977
rect 108684 291963 108712 296754
rect 109316 295384 109368 295390
rect 109316 295326 109368 295332
rect 109328 291963 109356 295326
rect 110340 294370 110368 340138
rect 110432 305794 110460 340711
rect 110420 305788 110472 305794
rect 110420 305730 110472 305736
rect 110524 303822 110552 378111
rect 110616 340785 110644 409838
rect 110696 387796 110748 387802
rect 110696 387738 110748 387744
rect 110708 353025 110736 387738
rect 111812 380934 111840 530538
rect 111984 396092 112036 396098
rect 111984 396034 112036 396040
rect 111892 391264 111944 391270
rect 111892 391206 111944 391212
rect 111800 380928 111852 380934
rect 111800 380870 111852 380876
rect 111798 378856 111854 378865
rect 111798 378791 111854 378800
rect 111812 378486 111840 378791
rect 111800 378480 111852 378486
rect 111800 378422 111852 378428
rect 111800 376848 111852 376854
rect 111798 376816 111800 376825
rect 111852 376816 111854 376825
rect 111798 376751 111854 376760
rect 111800 375760 111852 375766
rect 111800 375702 111852 375708
rect 111812 375465 111840 375702
rect 111798 375456 111854 375465
rect 111798 375391 111854 375400
rect 111798 374776 111854 374785
rect 111798 374711 111854 374720
rect 111812 374066 111840 374711
rect 111800 374060 111852 374066
rect 111800 374002 111852 374008
rect 111798 370016 111854 370025
rect 111798 369951 111800 369960
rect 111852 369951 111854 369960
rect 111800 369922 111852 369928
rect 111798 367296 111854 367305
rect 111798 367231 111854 367240
rect 111812 367130 111840 367231
rect 111800 367124 111852 367130
rect 111800 367066 111852 367072
rect 111798 365256 111854 365265
rect 111798 365191 111854 365200
rect 111812 364818 111840 365191
rect 111800 364812 111852 364818
rect 111800 364754 111852 364760
rect 111800 364676 111852 364682
rect 111800 364618 111852 364624
rect 110694 353016 110750 353025
rect 110694 352951 110750 352960
rect 111062 353016 111118 353025
rect 111062 352951 111118 352960
rect 111076 351966 111104 352951
rect 111064 351960 111116 351966
rect 111064 351902 111116 351908
rect 110602 340776 110658 340785
rect 110602 340711 110658 340720
rect 110512 303816 110564 303822
rect 110512 303758 110564 303764
rect 111708 303816 111760 303822
rect 111708 303758 111760 303764
rect 111720 301510 111748 303758
rect 111812 303006 111840 364618
rect 111904 364018 111932 391206
rect 111996 372842 112024 396034
rect 115204 392624 115256 392630
rect 115204 392566 115256 392572
rect 112444 389836 112496 389842
rect 112444 389778 112496 389784
rect 112168 380928 112220 380934
rect 112168 380870 112220 380876
rect 112074 376136 112130 376145
rect 112074 376071 112130 376080
rect 112088 375426 112116 376071
rect 112076 375420 112128 375426
rect 112076 375362 112128 375368
rect 112180 373994 112208 380870
rect 112088 373966 112208 373994
rect 111984 372836 112036 372842
rect 111984 372778 112036 372784
rect 111982 372736 112038 372745
rect 111982 372671 112038 372680
rect 111996 371226 112024 372671
rect 112088 371385 112116 373966
rect 112456 373425 112484 389778
rect 113916 387116 113968 387122
rect 113916 387058 113968 387064
rect 113824 382288 113876 382294
rect 113824 382230 113876 382236
rect 112442 373416 112498 373425
rect 112442 373351 112498 373360
rect 112168 372836 112220 372842
rect 112168 372778 112220 372784
rect 112074 371376 112130 371385
rect 112074 371311 112130 371320
rect 111996 371198 112116 371226
rect 111982 367976 112038 367985
rect 111982 367911 112038 367920
rect 111996 366353 112024 367911
rect 111982 366344 112038 366353
rect 111982 366279 112038 366288
rect 112088 364682 112116 371198
rect 112180 365945 112208 372778
rect 112352 372564 112404 372570
rect 112352 372506 112404 372512
rect 112364 372065 112392 372506
rect 112350 372056 112406 372065
rect 112350 371991 112406 372000
rect 112364 369170 112392 371991
rect 113086 370696 113142 370705
rect 113142 370654 113220 370682
rect 113086 370631 113142 370640
rect 112352 369164 112404 369170
rect 112352 369106 112404 369112
rect 112166 365936 112222 365945
rect 112166 365871 112222 365880
rect 112076 364676 112128 364682
rect 112076 364618 112128 364624
rect 111982 364576 112038 364585
rect 111982 364511 112038 364520
rect 111996 364410 112024 364511
rect 111984 364404 112036 364410
rect 111984 364346 112036 364352
rect 113192 364334 113220 370654
rect 113192 364306 113404 364334
rect 111904 363990 112208 364018
rect 112074 363896 112130 363905
rect 112074 363831 112130 363840
rect 111890 362536 111946 362545
rect 111890 362471 111946 362480
rect 111904 362302 111932 362471
rect 111892 362296 111944 362302
rect 111892 362238 111944 362244
rect 111984 362228 112036 362234
rect 111984 362170 112036 362176
rect 111996 361865 112024 362170
rect 111982 361856 112038 361865
rect 111982 361791 112038 361800
rect 111890 360496 111946 360505
rect 111890 360431 111946 360440
rect 111904 360330 111932 360431
rect 111892 360324 111944 360330
rect 111892 360266 111944 360272
rect 111982 359816 112038 359825
rect 111982 359751 112038 359760
rect 111890 359136 111946 359145
rect 111890 359071 111946 359080
rect 111904 358902 111932 359071
rect 111892 358896 111944 358902
rect 111892 358838 111944 358844
rect 111996 358834 112024 359751
rect 111984 358828 112036 358834
rect 111984 358770 112036 358776
rect 112088 358714 112116 363831
rect 111996 358686 112116 358714
rect 111892 357400 111944 357406
rect 111892 357342 111944 357348
rect 111904 357105 111932 357342
rect 111890 357096 111946 357105
rect 111890 357031 111946 357040
rect 111890 356416 111946 356425
rect 111890 356351 111946 356360
rect 111904 356114 111932 356351
rect 111892 356108 111944 356114
rect 111892 356050 111944 356056
rect 111890 355056 111946 355065
rect 111890 354991 111946 355000
rect 111904 354754 111932 354991
rect 111892 354748 111944 354754
rect 111892 354690 111944 354696
rect 111890 354376 111946 354385
rect 111890 354311 111946 354320
rect 111904 353326 111932 354311
rect 111892 353320 111944 353326
rect 111892 353262 111944 353268
rect 111890 351656 111946 351665
rect 111890 351591 111946 351600
rect 111904 350606 111932 351591
rect 111892 350600 111944 350606
rect 111892 350542 111944 350548
rect 111890 349616 111946 349625
rect 111890 349551 111946 349560
rect 111904 349178 111932 349551
rect 111892 349172 111944 349178
rect 111892 349114 111944 349120
rect 111890 348256 111946 348265
rect 111890 348191 111946 348200
rect 111904 347818 111932 348191
rect 111892 347812 111944 347818
rect 111892 347754 111944 347760
rect 111890 347576 111946 347585
rect 111890 347511 111946 347520
rect 111904 346458 111932 347511
rect 111892 346452 111944 346458
rect 111892 346394 111944 346400
rect 111890 345536 111946 345545
rect 111890 345471 111946 345480
rect 111904 345166 111932 345471
rect 111892 345160 111944 345166
rect 111892 345102 111944 345108
rect 111890 344856 111946 344865
rect 111890 344791 111946 344800
rect 111904 343874 111932 344791
rect 111996 344282 112024 358686
rect 112074 355736 112130 355745
rect 112074 355671 112130 355680
rect 111984 344276 112036 344282
rect 111984 344218 112036 344224
rect 111982 344176 112038 344185
rect 111982 344111 112038 344120
rect 111892 343868 111944 343874
rect 111892 343810 111944 343816
rect 111996 343670 112024 344111
rect 111984 343664 112036 343670
rect 111984 343606 112036 343612
rect 111892 343596 111944 343602
rect 111892 343538 111944 343544
rect 111904 343505 111932 343538
rect 111890 343496 111946 343505
rect 111890 343431 111946 343440
rect 111892 342236 111944 342242
rect 111892 342178 111944 342184
rect 111904 342145 111932 342178
rect 111890 342136 111946 342145
rect 111890 342071 111946 342080
rect 111890 340096 111946 340105
rect 111890 340031 111946 340040
rect 111904 303822 111932 340031
rect 112088 334762 112116 355671
rect 112180 354674 112208 363990
rect 112180 354646 112300 354674
rect 112166 350296 112222 350305
rect 112166 350231 112222 350240
rect 112180 349246 112208 350231
rect 112168 349240 112220 349246
rect 112168 349182 112220 349188
rect 112272 348945 112300 354646
rect 112258 348936 112314 348945
rect 112258 348871 112314 348880
rect 113270 348936 113326 348945
rect 113270 348871 113326 348880
rect 112166 346216 112222 346225
rect 112166 346151 112222 346160
rect 112180 345098 112208 346151
rect 112168 345092 112220 345098
rect 112168 345034 112220 345040
rect 112168 344276 112220 344282
rect 112168 344218 112220 344224
rect 112180 340202 112208 344218
rect 113086 342816 113142 342825
rect 113142 342774 113220 342802
rect 113086 342751 113142 342760
rect 112168 340196 112220 340202
rect 112168 340138 112220 340144
rect 113192 340105 113220 342774
rect 113178 340096 113234 340105
rect 113178 340031 113234 340040
rect 112076 334756 112128 334762
rect 112076 334698 112128 334704
rect 113284 330614 113312 348871
rect 113376 338842 113404 364306
rect 113836 358057 113864 382230
rect 113928 372570 113956 387058
rect 114652 379568 114704 379574
rect 114652 379510 114704 379516
rect 114008 378480 114060 378486
rect 114008 378422 114060 378428
rect 114020 373318 114048 378422
rect 114008 373312 114060 373318
rect 114008 373254 114060 373260
rect 113916 372564 113968 372570
rect 113916 372506 113968 372512
rect 114468 369980 114520 369986
rect 114468 369922 114520 369928
rect 114480 364993 114508 369922
rect 114466 364984 114522 364993
rect 114466 364919 114522 364928
rect 114560 364812 114612 364818
rect 114560 364754 114612 364760
rect 113822 358048 113878 358057
rect 113822 357983 113878 357992
rect 113364 338836 113416 338842
rect 113364 338778 113416 338784
rect 114572 337618 114600 364754
rect 114560 337612 114612 337618
rect 114560 337554 114612 337560
rect 113822 337376 113878 337385
rect 113822 337311 113878 337320
rect 113272 330608 113324 330614
rect 113272 330550 113324 330556
rect 113836 319433 113864 337311
rect 114560 324964 114612 324970
rect 114560 324906 114612 324912
rect 113822 319424 113878 319433
rect 113822 319359 113878 319368
rect 113824 308712 113876 308718
rect 113824 308654 113876 308660
rect 111892 303816 111944 303822
rect 111892 303758 111944 303764
rect 111800 303000 111852 303006
rect 111800 302942 111852 302948
rect 111708 301504 111760 301510
rect 111708 301446 111760 301452
rect 113836 298489 113864 308654
rect 113822 298480 113878 298489
rect 113822 298415 113878 298424
rect 111248 298308 111300 298314
rect 111248 298250 111300 298256
rect 110328 294364 110380 294370
rect 110328 294306 110380 294312
rect 110340 291977 110368 294306
rect 110604 292868 110656 292874
rect 110604 292810 110656 292816
rect 109986 291949 110368 291977
rect 110616 291963 110644 292810
rect 111260 291963 111288 298250
rect 111892 298240 111944 298246
rect 111892 298182 111944 298188
rect 111904 291963 111932 298182
rect 112536 296948 112588 296954
rect 112536 296890 112588 296896
rect 112548 291963 112576 296890
rect 113836 296714 113864 298415
rect 113744 296686 113864 296714
rect 113744 291977 113772 296686
rect 114468 294228 114520 294234
rect 114468 294170 114520 294176
rect 114376 294024 114428 294030
rect 114376 293966 114428 293972
rect 113206 291949 113772 291977
rect 114388 291977 114416 293966
rect 114480 293282 114508 294170
rect 114468 293276 114520 293282
rect 114468 293218 114520 293224
rect 114572 291977 114600 324906
rect 114664 296818 114692 379510
rect 115216 338094 115244 392566
rect 115860 383654 115888 702578
rect 116584 470620 116636 470626
rect 116584 470562 116636 470568
rect 115768 383626 115888 383654
rect 115294 382392 115350 382401
rect 115294 382327 115350 382336
rect 115308 352617 115336 382327
rect 115768 376786 115796 383626
rect 115756 376780 115808 376786
rect 115756 376722 115808 376728
rect 115768 375766 115796 376722
rect 115756 375760 115808 375766
rect 115756 375702 115808 375708
rect 116596 362234 116624 470562
rect 116676 375420 116728 375426
rect 116676 375362 116728 375368
rect 116584 362228 116636 362234
rect 116584 362170 116636 362176
rect 115294 352608 115350 352617
rect 115294 352543 115350 352552
rect 115848 343868 115900 343874
rect 115848 343810 115900 343816
rect 115860 342922 115888 343810
rect 115848 342916 115900 342922
rect 115848 342858 115900 342864
rect 115204 338088 115256 338094
rect 115204 338030 115256 338036
rect 115204 329248 115256 329254
rect 115204 329190 115256 329196
rect 115216 306374 115244 329190
rect 115940 312588 115992 312594
rect 115940 312530 115992 312536
rect 115216 306346 115336 306374
rect 114652 296812 114704 296818
rect 114652 296754 114704 296760
rect 115308 294273 115336 306346
rect 115294 294264 115350 294273
rect 115294 294199 115350 294208
rect 114190 291952 114246 291961
rect 79336 291910 79706 291938
rect 80624 291910 80994 291938
rect 81912 291910 82282 291938
rect 84304 291910 84858 291938
rect 85592 291910 86146 291938
rect 94792 291910 95162 291938
rect 97368 291910 97738 291938
rect 102336 291910 102890 291938
rect 103624 291910 104178 291938
rect 106384 291910 106754 291938
rect 108304 291916 108356 291922
rect 108054 291864 108304 291870
rect 113850 291910 114190 291938
rect 114388 291949 114494 291977
rect 114572 291949 115138 291977
rect 115308 291938 115336 294199
rect 115952 291977 115980 312530
rect 116596 293457 116624 362170
rect 116688 303822 116716 375362
rect 117240 342242 117268 702850
rect 123484 702772 123536 702778
rect 123484 702714 123536 702720
rect 119988 702704 120040 702710
rect 119988 702646 120040 702652
rect 118608 391264 118660 391270
rect 118608 391206 118660 391212
rect 117320 388476 117372 388482
rect 117320 388418 117372 388424
rect 117228 342236 117280 342242
rect 117228 342178 117280 342184
rect 117240 340950 117268 342178
rect 117228 340944 117280 340950
rect 117228 340886 117280 340892
rect 117332 339318 117360 388418
rect 118620 373994 118648 391206
rect 118700 383852 118752 383858
rect 118700 383794 118752 383800
rect 118528 373966 118648 373994
rect 118528 357474 118556 373966
rect 118608 365764 118660 365770
rect 118608 365706 118660 365712
rect 118620 362234 118648 365706
rect 118608 362228 118660 362234
rect 118608 362170 118660 362176
rect 118516 357468 118568 357474
rect 118516 357410 118568 357416
rect 117320 339312 117372 339318
rect 117320 339254 117372 339260
rect 118712 306374 118740 383794
rect 119344 376848 119396 376854
rect 119344 376790 119396 376796
rect 119356 363662 119384 376790
rect 119344 363656 119396 363662
rect 119344 363598 119396 363604
rect 120000 343777 120028 702646
rect 122104 536852 122156 536858
rect 122104 536794 122156 536800
rect 121460 385348 121512 385354
rect 121460 385290 121512 385296
rect 120080 369164 120132 369170
rect 120080 369106 120132 369112
rect 119986 343768 120042 343777
rect 119986 343703 120042 343712
rect 120000 343602 120028 343703
rect 119988 343596 120040 343602
rect 119988 343538 120040 343544
rect 118712 306346 119200 306374
rect 117412 305720 117464 305726
rect 117412 305662 117464 305668
rect 116676 303816 116728 303822
rect 116676 303758 116728 303764
rect 117320 303816 117372 303822
rect 117320 303758 117372 303764
rect 117044 296812 117096 296818
rect 117044 296754 117096 296760
rect 116582 293448 116638 293457
rect 116582 293383 116638 293392
rect 115952 291949 116426 291977
rect 117056 291963 117084 296754
rect 117332 295662 117360 303758
rect 117424 298110 117452 305662
rect 117412 298104 117464 298110
rect 117412 298046 117464 298052
rect 117320 295656 117372 295662
rect 117320 295598 117372 295604
rect 118332 295656 118384 295662
rect 118332 295598 118384 295604
rect 117964 294432 118016 294438
rect 117964 294374 118016 294380
rect 117688 292800 117740 292806
rect 117688 292742 117740 292748
rect 117700 291963 117728 292742
rect 115308 291910 115770 291938
rect 117976 291922 118004 294374
rect 118344 291963 118372 295598
rect 118976 294228 119028 294234
rect 118976 294170 119028 294176
rect 118988 291963 119016 294170
rect 119172 291938 119200 306346
rect 119804 294364 119856 294370
rect 119804 294306 119856 294312
rect 117964 291916 118016 291922
rect 114190 291887 114246 291896
rect 108054 291858 108356 291864
rect 119172 291910 119646 291938
rect 117964 291858 118016 291864
rect 108054 291842 108344 291858
rect 69018 291136 69074 291145
rect 69018 291071 69074 291080
rect 119816 289134 119844 294306
rect 119804 289128 119856 289134
rect 119804 289070 119856 289076
rect 68742 286104 68798 286113
rect 68742 286039 68798 286048
rect 68650 284744 68706 284753
rect 68650 284679 68706 284688
rect 67640 284300 67692 284306
rect 67640 284242 67692 284248
rect 67652 283393 67680 284242
rect 68926 283792 68982 283801
rect 68926 283727 68982 283736
rect 67638 283384 67694 283393
rect 67638 283319 67694 283328
rect 67640 282872 67692 282878
rect 67640 282814 67692 282820
rect 67652 282169 67680 282814
rect 67638 282160 67694 282169
rect 67638 282095 67694 282104
rect 68282 280528 68338 280537
rect 68282 280463 68338 280472
rect 67638 280392 67694 280401
rect 67638 280327 67694 280336
rect 67652 280226 67680 280327
rect 67640 280220 67692 280226
rect 67640 280162 67692 280168
rect 67732 280152 67784 280158
rect 67732 280094 67784 280100
rect 67640 280084 67692 280090
rect 67640 280026 67692 280032
rect 67652 279313 67680 280026
rect 67744 279993 67772 280094
rect 67730 279984 67786 279993
rect 67730 279919 67786 279928
rect 67638 279304 67694 279313
rect 67638 279239 67694 279248
rect 67730 277808 67786 277817
rect 67730 277743 67786 277752
rect 67638 277672 67694 277681
rect 67638 277607 67694 277616
rect 67652 277506 67680 277607
rect 67640 277500 67692 277506
rect 67640 277442 67692 277448
rect 67744 277438 67772 277743
rect 67732 277432 67784 277438
rect 67732 277374 67784 277380
rect 67638 276448 67694 276457
rect 67638 276383 67694 276392
rect 67652 276146 67680 276383
rect 67640 276140 67692 276146
rect 67640 276082 67692 276088
rect 67822 275088 67878 275097
rect 67822 275023 67878 275032
rect 67638 274952 67694 274961
rect 67638 274887 67694 274896
rect 67652 274786 67680 274887
rect 67640 274780 67692 274786
rect 67640 274722 67692 274728
rect 67836 274718 67864 275023
rect 67824 274712 67876 274718
rect 67824 274654 67876 274660
rect 67732 274644 67784 274650
rect 67732 274586 67784 274592
rect 67744 274553 67772 274586
rect 67730 274544 67786 274553
rect 67730 274479 67786 274488
rect 67822 272368 67878 272377
rect 67822 272303 67878 272312
rect 67638 272232 67694 272241
rect 67638 272167 67694 272176
rect 67652 271998 67680 272167
rect 67640 271992 67692 271998
rect 67640 271934 67692 271940
rect 67836 271930 67864 272303
rect 67824 271924 67876 271930
rect 67824 271866 67876 271872
rect 67732 271856 67784 271862
rect 67732 271798 67784 271804
rect 67638 271008 67694 271017
rect 67638 270943 67694 270952
rect 67652 270570 67680 270943
rect 67744 270881 67772 271798
rect 67730 270872 67786 270881
rect 67730 270807 67786 270816
rect 67640 270564 67692 270570
rect 67640 270506 67692 270512
rect 67730 269648 67786 269657
rect 67730 269583 67786 269592
rect 67638 269512 67694 269521
rect 67638 269447 67694 269456
rect 67652 269142 67680 269447
rect 67744 269210 67772 269583
rect 67732 269204 67784 269210
rect 67732 269146 67784 269152
rect 67640 269136 67692 269142
rect 67640 269078 67692 269084
rect 67640 268388 67692 268394
rect 67640 268330 67692 268336
rect 67652 268161 67680 268330
rect 68190 268288 68246 268297
rect 68190 268223 68192 268232
rect 68244 268223 68246 268232
rect 68192 268194 68244 268200
rect 67638 268152 67694 268161
rect 67638 268087 67694 268096
rect 67732 267708 67784 267714
rect 67732 267650 67784 267656
rect 67640 267640 67692 267646
rect 67638 267608 67640 267617
rect 67692 267608 67694 267617
rect 67638 267543 67694 267552
rect 67744 267073 67772 267650
rect 67730 267064 67786 267073
rect 67730 266999 67786 267008
rect 67640 266348 67692 266354
rect 67640 266290 67692 266296
rect 67652 265441 67680 266290
rect 67730 265568 67786 265577
rect 67730 265503 67786 265512
rect 67638 265432 67694 265441
rect 67638 265367 67694 265376
rect 67744 264994 67772 265503
rect 67732 264988 67784 264994
rect 67732 264930 67784 264936
rect 67640 264920 67692 264926
rect 67638 264888 67640 264897
rect 67692 264888 67694 264897
rect 67638 264823 67694 264832
rect 67730 263664 67786 263673
rect 67730 263599 67732 263608
rect 67784 263599 67786 263608
rect 67732 263570 67784 263576
rect 67640 263560 67692 263566
rect 67638 263528 67640 263537
rect 67692 263528 67694 263537
rect 67638 263463 67694 263472
rect 67638 262304 67694 262313
rect 67638 262239 67640 262248
rect 67692 262239 67694 262248
rect 67640 262210 67692 262216
rect 67638 261488 67694 261497
rect 67638 261423 67694 261432
rect 67652 260982 67680 261423
rect 67640 260976 67692 260982
rect 67640 260918 67692 260924
rect 67730 260944 67786 260953
rect 67730 260879 67732 260888
rect 67784 260879 67786 260888
rect 67732 260850 67784 260856
rect 67640 260840 67692 260846
rect 67638 260808 67640 260817
rect 67692 260808 67694 260817
rect 67638 260743 67694 260752
rect 67638 259584 67694 259593
rect 67638 259519 67694 259528
rect 67652 259486 67680 259519
rect 67640 259480 67692 259486
rect 67640 259422 67692 259428
rect 67730 258632 67786 258641
rect 67730 258567 67786 258576
rect 67638 258224 67694 258233
rect 67638 258159 67640 258168
rect 67692 258159 67694 258168
rect 67640 258130 67692 258136
rect 67744 258126 67772 258567
rect 67732 258120 67784 258126
rect 67732 258062 67784 258068
rect 67640 258052 67692 258058
rect 67640 257994 67692 258000
rect 67652 257961 67680 257994
rect 67638 257952 67694 257961
rect 67638 257887 67694 257896
rect 68296 257378 68324 280463
rect 68374 273592 68430 273601
rect 68374 273527 68430 273536
rect 68388 257446 68416 273527
rect 68376 257440 68428 257446
rect 68376 257382 68428 257388
rect 68284 257372 68336 257378
rect 68284 257314 68336 257320
rect 67638 256864 67694 256873
rect 67638 256799 67694 256808
rect 67652 256766 67680 256799
rect 67640 256760 67692 256766
rect 67640 256702 67692 256708
rect 68834 255368 68890 255377
rect 68834 255303 68890 255312
rect 67640 255264 67692 255270
rect 67638 255232 67640 255241
rect 67692 255232 67694 255241
rect 67638 255167 67694 255176
rect 67640 254652 67692 254658
rect 67640 254594 67692 254600
rect 67652 254561 67680 254594
rect 67638 254552 67694 254561
rect 67638 254487 67694 254496
rect 67640 253904 67692 253910
rect 67638 253872 67640 253881
rect 67692 253872 67694 253881
rect 67638 253807 67694 253816
rect 67638 252648 67694 252657
rect 67638 252583 67640 252592
rect 67692 252583 67694 252592
rect 67640 252554 67692 252560
rect 67730 251832 67786 251841
rect 67730 251767 67786 251776
rect 67744 251326 67772 251767
rect 67732 251320 67784 251326
rect 67638 251288 67694 251297
rect 67732 251262 67784 251268
rect 67638 251223 67640 251232
rect 67692 251223 67694 251232
rect 67640 251194 67692 251200
rect 67638 250472 67694 250481
rect 67638 250407 67694 250416
rect 67652 249898 67680 250407
rect 67730 249928 67786 249937
rect 67640 249892 67692 249898
rect 67730 249863 67786 249872
rect 67640 249834 67692 249840
rect 67744 249830 67772 249863
rect 67732 249824 67784 249830
rect 67638 249792 67694 249801
rect 67732 249766 67784 249772
rect 67638 249727 67640 249736
rect 67692 249727 67694 249736
rect 67640 249698 67692 249704
rect 68098 248704 68154 248713
rect 68098 248639 68100 248648
rect 68152 248639 68154 248648
rect 68100 248610 68152 248616
rect 67730 247752 67786 247761
rect 67730 247687 67786 247696
rect 67638 247208 67694 247217
rect 67744 247178 67772 247687
rect 67638 247143 67694 247152
rect 67732 247172 67784 247178
rect 67652 247110 67680 247143
rect 67732 247114 67784 247120
rect 67640 247104 67692 247110
rect 67640 247046 67692 247052
rect 67640 245608 67692 245614
rect 67640 245550 67692 245556
rect 67652 245313 67680 245550
rect 67638 245304 67694 245313
rect 67638 245239 67694 245248
rect 68098 244352 68154 244361
rect 68098 244287 68100 244296
rect 68152 244287 68154 244296
rect 68100 244258 68152 244264
rect 67640 244248 67692 244254
rect 67640 244190 67692 244196
rect 67652 243273 67680 244190
rect 67638 243264 67694 243273
rect 67638 243199 67694 243208
rect 67638 241904 67694 241913
rect 67638 241839 67694 241848
rect 67652 241534 67680 241839
rect 67640 241528 67692 241534
rect 67640 241470 67692 241476
rect 68848 238066 68876 255303
rect 68836 238060 68888 238066
rect 68836 238002 68888 238008
rect 68940 236706 68968 283727
rect 69018 255912 69074 255921
rect 69018 255847 69074 255856
rect 68928 236700 68980 236706
rect 68928 236642 68980 236648
rect 69032 196722 69060 255847
rect 120092 252385 120120 369106
rect 120724 340944 120776 340950
rect 120724 340886 120776 340892
rect 120170 293312 120226 293321
rect 120170 293247 120226 293256
rect 120184 285705 120212 293247
rect 120170 285696 120226 285705
rect 120170 285631 120226 285640
rect 120078 252376 120134 252385
rect 120078 252311 120134 252320
rect 120448 251048 120500 251054
rect 120078 251016 120134 251025
rect 120078 250951 120134 250960
rect 120446 251016 120448 251025
rect 120500 251016 120502 251025
rect 120446 250951 120502 250960
rect 69110 245712 69166 245721
rect 69110 245647 69166 245656
rect 69020 196716 69072 196722
rect 69020 196658 69072 196664
rect 69124 188426 69152 245647
rect 69202 243672 69258 243681
rect 69202 243607 69258 243616
rect 69216 188494 69244 243607
rect 69754 240272 69810 240281
rect 69754 240207 69810 240216
rect 69768 239562 69796 240207
rect 119896 240168 119948 240174
rect 69952 240094 70058 240122
rect 119646 240116 119896 240122
rect 119646 240110 119948 240116
rect 119646 240094 119936 240110
rect 69756 239556 69808 239562
rect 69756 239498 69808 239504
rect 69952 237454 69980 240094
rect 70688 238754 70716 240037
rect 70412 238726 70716 238754
rect 69940 237448 69992 237454
rect 69940 237390 69992 237396
rect 70412 192506 70440 238726
rect 71332 237522 71360 240037
rect 71964 239850 71992 240037
rect 72516 239964 72568 239970
rect 72516 239906 72568 239912
rect 71884 239822 71992 239850
rect 71320 237516 71372 237522
rect 71320 237458 71372 237464
rect 70400 192500 70452 192506
rect 70400 192442 70452 192448
rect 69204 188488 69256 188494
rect 69204 188430 69256 188436
rect 69112 188420 69164 188426
rect 69112 188362 69164 188368
rect 67548 184340 67600 184346
rect 67548 184282 67600 184288
rect 71884 180130 71912 239822
rect 72424 237448 72476 237454
rect 72424 237390 72476 237396
rect 72436 202162 72464 237390
rect 72528 229770 72556 239906
rect 72620 238610 72648 240037
rect 73252 239850 73280 240037
rect 73896 239850 73924 240037
rect 73172 239822 73280 239850
rect 73816 239822 73924 239850
rect 72608 238604 72660 238610
rect 72608 238546 72660 238552
rect 72516 229764 72568 229770
rect 72516 229706 72568 229712
rect 72424 202156 72476 202162
rect 72424 202098 72476 202104
rect 73172 184278 73200 239822
rect 73816 219434 73844 239822
rect 73264 219406 73844 219434
rect 73264 186998 73292 219406
rect 73252 186992 73304 186998
rect 73252 186934 73304 186940
rect 73160 184272 73212 184278
rect 73160 184214 73212 184220
rect 74552 181393 74580 240037
rect 75196 238754 75224 240037
rect 74644 238726 75224 238754
rect 74644 207670 74672 238726
rect 75184 237516 75236 237522
rect 75184 237458 75236 237464
rect 75196 221542 75224 237458
rect 75840 237386 75868 240037
rect 75920 239828 75972 239834
rect 75920 239770 75972 239776
rect 75828 237380 75880 237386
rect 75828 237322 75880 237328
rect 75184 221536 75236 221542
rect 75184 221478 75236 221484
rect 74632 207664 74684 207670
rect 74632 207606 74684 207612
rect 75932 182850 75960 239770
rect 76484 238754 76512 240037
rect 77116 239834 77144 240037
rect 77104 239828 77156 239834
rect 77104 239770 77156 239776
rect 77772 238754 77800 240037
rect 78404 239816 78432 240037
rect 76484 238726 76604 238754
rect 76576 235754 76604 238726
rect 77312 238726 77800 238754
rect 78324 239788 78432 239816
rect 78680 239828 78732 239834
rect 76564 235748 76616 235754
rect 76564 235690 76616 235696
rect 76576 198014 76604 235690
rect 77312 199442 77340 238726
rect 78324 231130 78352 239788
rect 78680 239770 78732 239776
rect 78312 231124 78364 231130
rect 78312 231066 78364 231072
rect 77300 199436 77352 199442
rect 77300 199378 77352 199384
rect 76564 198008 76616 198014
rect 76564 197950 76616 197956
rect 78692 193866 78720 239770
rect 79060 238754 79088 240037
rect 79692 239834 79720 240037
rect 79680 239828 79732 239834
rect 79680 239770 79732 239776
rect 78784 238726 79088 238754
rect 78784 224330 78812 238726
rect 80348 233986 80376 240037
rect 80980 239816 81008 240037
rect 80900 239788 81008 239816
rect 80336 233980 80388 233986
rect 80336 233922 80388 233928
rect 78772 224324 78824 224330
rect 78772 224266 78824 224272
rect 80900 219434 80928 239788
rect 81636 235754 81664 240037
rect 82082 239456 82138 239465
rect 82082 239391 82138 239400
rect 81624 235748 81676 235754
rect 81624 235690 81676 235696
rect 80072 219406 80928 219434
rect 78680 193860 78732 193866
rect 78680 193802 78732 193808
rect 80072 185706 80100 219406
rect 82096 217326 82124 239391
rect 82280 238678 82308 240037
rect 82268 238672 82320 238678
rect 82268 238614 82320 238620
rect 82924 238134 82952 240037
rect 83568 239714 83596 240037
rect 83476 239686 83596 239714
rect 83476 238754 83504 239686
rect 83556 239556 83608 239562
rect 83556 239498 83608 239504
rect 83384 238726 83504 238754
rect 82912 238128 82964 238134
rect 82912 238070 82964 238076
rect 83384 230450 83412 238726
rect 83372 230444 83424 230450
rect 83372 230386 83424 230392
rect 83568 219434 83596 239498
rect 84212 239442 84240 240037
rect 84212 239414 84424 239442
rect 84292 239352 84344 239358
rect 84292 239294 84344 239300
rect 84108 231872 84160 231878
rect 84160 231826 84240 231854
rect 84108 231814 84160 231820
rect 83476 219406 83596 219434
rect 82084 217320 82136 217326
rect 82084 217262 82136 217268
rect 83476 210458 83504 219406
rect 83464 210452 83516 210458
rect 83464 210394 83516 210400
rect 80060 185700 80112 185706
rect 80060 185642 80112 185648
rect 84212 182918 84240 231826
rect 84304 192574 84332 239294
rect 84396 226953 84424 239414
rect 84856 231878 84884 240037
rect 85500 239358 85528 240037
rect 85488 239352 85540 239358
rect 85488 239294 85540 239300
rect 86144 238754 86172 240037
rect 86144 238726 86264 238754
rect 86788 238746 86816 240037
rect 86960 239828 87012 239834
rect 86960 239770 87012 239776
rect 86236 237289 86264 238726
rect 86776 238740 86828 238746
rect 86776 238682 86828 238688
rect 86222 237280 86278 237289
rect 86222 237215 86278 237224
rect 84844 231872 84896 231878
rect 84844 231814 84896 231820
rect 84382 226944 84438 226953
rect 84382 226879 84438 226888
rect 86236 195294 86264 237215
rect 86972 207738 87000 239770
rect 87432 238754 87460 240037
rect 88064 239834 88092 240037
rect 88052 239828 88104 239834
rect 88052 239770 88104 239776
rect 88720 238754 88748 240037
rect 87064 238726 87460 238754
rect 88352 238726 88748 238754
rect 89364 238746 89392 240037
rect 89720 239828 89772 239834
rect 89720 239770 89772 239776
rect 89352 238740 89404 238746
rect 87064 213314 87092 238726
rect 88352 228410 88380 238726
rect 89352 238682 89404 238688
rect 88984 238128 89036 238134
rect 88984 238070 89036 238076
rect 88996 234530 89024 238070
rect 88984 234524 89036 234530
rect 88984 234466 89036 234472
rect 88340 228404 88392 228410
rect 88340 228346 88392 228352
rect 87052 213308 87104 213314
rect 87052 213250 87104 213256
rect 86960 207732 87012 207738
rect 86960 207674 87012 207680
rect 89732 205018 89760 239770
rect 90008 238754 90036 240037
rect 90640 239834 90668 240037
rect 90628 239828 90680 239834
rect 90628 239770 90680 239776
rect 89824 238726 90036 238754
rect 89824 213382 89852 238726
rect 91296 235686 91324 240037
rect 91940 238678 91968 240037
rect 92572 239850 92600 240037
rect 93216 239850 93244 240037
rect 92492 239822 92600 239850
rect 93136 239822 93244 239850
rect 91928 238672 91980 238678
rect 91928 238614 91980 238620
rect 91940 238513 91968 238614
rect 91926 238504 91982 238513
rect 91926 238439 91982 238448
rect 91284 235680 91336 235686
rect 91284 235622 91336 235628
rect 89812 213376 89864 213382
rect 89812 213318 89864 213324
rect 89720 205012 89772 205018
rect 89720 204954 89772 204960
rect 92492 196790 92520 239822
rect 93136 219434 93164 239822
rect 92584 219406 93164 219434
rect 92584 198082 92612 219406
rect 93872 200938 93900 240037
rect 94516 238754 94544 240037
rect 95148 239816 95176 240037
rect 93964 238726 94544 238754
rect 95068 239788 95176 239816
rect 93964 215966 93992 238726
rect 95068 224262 95096 239788
rect 95804 238814 95832 240037
rect 95792 238808 95844 238814
rect 95792 238750 95844 238756
rect 96448 238134 96476 240037
rect 97092 238754 97120 240037
rect 97724 239816 97752 240037
rect 96632 238726 97120 238754
rect 97644 239788 97752 239816
rect 96436 238128 96488 238134
rect 96436 238070 96488 238076
rect 95056 224256 95108 224262
rect 95056 224198 95108 224204
rect 93952 215960 94004 215966
rect 93952 215902 94004 215908
rect 93860 200932 93912 200938
rect 93860 200874 93912 200880
rect 96632 200870 96660 238726
rect 97644 228478 97672 239788
rect 98380 238649 98408 240037
rect 99024 239018 99052 240037
rect 99012 239012 99064 239018
rect 99012 238954 99064 238960
rect 99668 238754 99696 240037
rect 100300 239816 100328 240037
rect 99392 238726 99696 238754
rect 100220 239788 100328 239816
rect 100760 239828 100812 239834
rect 98366 238640 98422 238649
rect 98366 238575 98422 238584
rect 97632 228472 97684 228478
rect 97632 228414 97684 228420
rect 96620 200864 96672 200870
rect 96620 200806 96672 200812
rect 92572 198076 92624 198082
rect 92572 198018 92624 198024
rect 92480 196784 92532 196790
rect 92480 196726 92532 196732
rect 86224 195288 86276 195294
rect 86224 195230 86276 195236
rect 84292 192568 84344 192574
rect 84292 192510 84344 192516
rect 99288 186448 99340 186454
rect 99288 186390 99340 186396
rect 84200 182912 84252 182918
rect 84200 182854 84252 182860
rect 75920 182844 75972 182850
rect 75920 182786 75972 182792
rect 74538 181384 74594 181393
rect 74538 181319 74594 181328
rect 71872 180124 71924 180130
rect 71872 180066 71924 180072
rect 97262 179480 97318 179489
rect 97262 179415 97318 179424
rect 66168 178764 66220 178770
rect 66168 178706 66220 178712
rect 97276 177041 97304 179415
rect 99300 177721 99328 186390
rect 99392 185842 99420 238726
rect 100220 219434 100248 239788
rect 100944 239816 100972 240037
rect 101588 239834 101616 240037
rect 100760 239770 100812 239776
rect 100864 239788 100972 239816
rect 101576 239828 101628 239834
rect 99484 219406 100248 219434
rect 99484 216034 99512 219406
rect 99472 216028 99524 216034
rect 99472 215970 99524 215976
rect 100772 202230 100800 239770
rect 100864 209234 100892 239788
rect 102232 239816 102260 240037
rect 101576 239770 101628 239776
rect 102152 239788 102260 239816
rect 100852 209228 100904 209234
rect 100852 209170 100904 209176
rect 100760 202224 100812 202230
rect 100760 202166 100812 202172
rect 100668 186516 100720 186522
rect 100668 186458 100720 186464
rect 99380 185836 99432 185842
rect 99380 185778 99432 185784
rect 99286 177712 99342 177721
rect 99286 177647 99342 177656
rect 97262 177032 97318 177041
rect 97262 176967 97318 176976
rect 100680 176769 100708 186458
rect 102152 178702 102180 239788
rect 102888 238202 102916 240037
rect 102876 238196 102928 238202
rect 102876 238138 102928 238144
rect 103532 235958 103560 240037
rect 103612 239828 103664 239834
rect 103612 239770 103664 239776
rect 103520 235952 103572 235958
rect 103520 235894 103572 235900
rect 103624 218754 103652 239770
rect 104176 238754 104204 240037
rect 104808 239834 104836 240037
rect 104796 239828 104848 239834
rect 104796 239770 104848 239776
rect 104900 239828 104952 239834
rect 104900 239770 104952 239776
rect 103716 238726 104204 238754
rect 103612 218748 103664 218754
rect 103612 218690 103664 218696
rect 103716 214606 103744 238726
rect 103704 214600 103756 214606
rect 103704 214542 103756 214548
rect 104808 187740 104860 187746
rect 104808 187682 104860 187688
rect 102140 178696 102192 178702
rect 102140 178638 102192 178644
rect 104820 177721 104848 187682
rect 104912 185774 104940 239770
rect 105464 238754 105492 240037
rect 106096 239834 106124 240037
rect 106084 239828 106136 239834
rect 106084 239770 106136 239776
rect 105004 238726 105492 238754
rect 105004 211818 105032 238726
rect 106752 238542 106780 240037
rect 106740 238536 106792 238542
rect 106740 238478 106792 238484
rect 106924 238196 106976 238202
rect 106924 238138 106976 238144
rect 104992 211812 105044 211818
rect 104992 211754 105044 211760
rect 106936 202298 106964 238138
rect 107396 235822 107424 240037
rect 107660 239828 107712 239834
rect 107660 239770 107712 239776
rect 107384 235816 107436 235822
rect 107384 235758 107436 235764
rect 106924 202292 106976 202298
rect 106924 202234 106976 202240
rect 107672 196654 107700 239770
rect 108040 238754 108068 240037
rect 108672 239834 108700 240037
rect 108660 239828 108712 239834
rect 108660 239770 108712 239776
rect 107764 238726 108068 238754
rect 107764 200802 107792 238726
rect 109040 234592 109092 234598
rect 109040 234534 109092 234540
rect 109052 234190 109080 234534
rect 109972 234190 110000 240037
rect 110616 234598 110644 240037
rect 111260 238754 111288 240037
rect 111892 239850 111920 240037
rect 110892 238726 111288 238754
rect 111812 239822 111920 239850
rect 110604 234592 110656 234598
rect 110604 234534 110656 234540
rect 109040 234184 109092 234190
rect 109040 234126 109092 234132
rect 109960 234184 110012 234190
rect 109960 234126 110012 234132
rect 107752 200796 107804 200802
rect 107752 200738 107804 200744
rect 107660 196648 107712 196654
rect 107660 196590 107712 196596
rect 107568 189100 107620 189106
rect 107568 189042 107620 189048
rect 104900 185768 104952 185774
rect 104900 185710 104952 185716
rect 107580 177721 107608 189042
rect 109052 188562 109080 234126
rect 110892 219434 110920 238726
rect 111064 234592 111116 234598
rect 111064 234534 111116 234540
rect 110432 219406 110920 219434
rect 110432 218822 110460 219406
rect 110420 218816 110472 218822
rect 110420 218758 110472 218764
rect 109040 188556 109092 188562
rect 109040 188498 109092 188504
rect 110696 182232 110748 182238
rect 110696 182174 110748 182180
rect 110052 178084 110104 178090
rect 110052 178026 110104 178032
rect 104806 177712 104862 177721
rect 104806 177647 104862 177656
rect 107566 177712 107622 177721
rect 107566 177647 107622 177656
rect 103336 176996 103388 177002
rect 103336 176938 103388 176944
rect 103348 176769 103376 176938
rect 108120 176928 108172 176934
rect 108120 176870 108172 176876
rect 108132 176769 108160 176870
rect 110064 176769 110092 178026
rect 110708 177721 110736 182174
rect 110694 177712 110750 177721
rect 110694 177647 110750 177656
rect 100666 176760 100722 176769
rect 100666 176695 100722 176704
rect 102046 176760 102102 176769
rect 102046 176695 102048 176704
rect 102100 176695 102102 176704
rect 103334 176760 103390 176769
rect 103334 176695 103390 176704
rect 108118 176760 108174 176769
rect 108118 176695 108174 176704
rect 110050 176760 110106 176769
rect 110050 176695 110106 176704
rect 102048 176666 102100 176672
rect 100760 176044 100812 176050
rect 100760 175986 100812 175992
rect 100772 175409 100800 175986
rect 111076 175982 111104 234534
rect 111812 206310 111840 239822
rect 112548 235890 112576 240037
rect 112536 235884 112588 235890
rect 112536 235826 112588 235832
rect 113192 209098 113220 240037
rect 113836 238649 113864 240037
rect 114480 238882 114508 240037
rect 114560 239828 114612 239834
rect 114560 239770 114612 239776
rect 114468 238876 114520 238882
rect 114468 238818 114520 238824
rect 113822 238640 113878 238649
rect 113822 238575 113878 238584
rect 114572 220182 114600 239770
rect 115124 238950 115152 240037
rect 115756 239834 115784 240037
rect 115744 239828 115796 239834
rect 115744 239770 115796 239776
rect 115112 238944 115164 238950
rect 115112 238886 115164 238892
rect 116412 238754 116440 240037
rect 115952 238726 116440 238754
rect 114560 220176 114612 220182
rect 114560 220118 114612 220124
rect 113180 209092 113232 209098
rect 113180 209034 113232 209040
rect 111800 206304 111852 206310
rect 111800 206246 111852 206252
rect 115952 199510 115980 238726
rect 117056 238513 117084 240037
rect 117042 238504 117098 238513
rect 117042 238439 117098 238448
rect 117700 235958 117728 240037
rect 118344 238610 118372 240037
rect 118976 239873 119004 240037
rect 118962 239864 119018 239873
rect 118962 239799 119018 239808
rect 118332 238604 118384 238610
rect 118332 238546 118384 238552
rect 117688 235952 117740 235958
rect 117688 235894 117740 235900
rect 120092 225622 120120 250951
rect 120736 249558 120764 340886
rect 121472 308446 121500 385290
rect 121552 379636 121604 379642
rect 121552 379578 121604 379584
rect 121564 323746 121592 379578
rect 122116 362302 122144 536794
rect 122840 380996 122892 381002
rect 122840 380938 122892 380944
rect 122104 362296 122156 362302
rect 122104 362238 122156 362244
rect 121552 323740 121604 323746
rect 121552 323682 121604 323688
rect 121828 323740 121880 323746
rect 121828 323682 121880 323688
rect 121840 323610 121868 323682
rect 121828 323604 121880 323610
rect 121828 323546 121880 323552
rect 121644 309868 121696 309874
rect 121644 309810 121696 309816
rect 121460 308440 121512 308446
rect 121460 308382 121512 308388
rect 121552 298104 121604 298110
rect 121552 298046 121604 298052
rect 121460 292528 121512 292534
rect 121460 292470 121512 292476
rect 121472 291825 121500 292470
rect 121458 291816 121514 291825
rect 121458 291751 121514 291760
rect 121458 291136 121514 291145
rect 121458 291071 121514 291080
rect 121472 289950 121500 291071
rect 121460 289944 121512 289950
rect 121460 289886 121512 289892
rect 121460 289808 121512 289814
rect 121458 289776 121460 289785
rect 121512 289776 121514 289785
rect 121458 289711 121514 289720
rect 121460 288380 121512 288386
rect 121460 288322 121512 288328
rect 121472 287745 121500 288322
rect 121458 287736 121514 287745
rect 121458 287671 121514 287680
rect 121458 287056 121514 287065
rect 121458 286991 121460 287000
rect 121512 286991 121514 287000
rect 121460 286962 121512 286968
rect 120908 286408 120960 286414
rect 121564 286385 121592 298046
rect 120908 286350 120960 286356
rect 121550 286376 121606 286385
rect 120816 285728 120868 285734
rect 120814 285696 120816 285705
rect 120868 285696 120870 285705
rect 120814 285631 120870 285640
rect 120920 277394 120948 286350
rect 121550 286311 121606 286320
rect 121550 285016 121606 285025
rect 121550 284951 121606 284960
rect 121564 284374 121592 284951
rect 121552 284368 121604 284374
rect 121552 284310 121604 284316
rect 121460 284300 121512 284306
rect 121460 284242 121512 284248
rect 121472 283665 121500 284242
rect 121458 283656 121514 283665
rect 121458 283591 121514 283600
rect 121458 282976 121514 282985
rect 121458 282911 121460 282920
rect 121512 282911 121514 282920
rect 121460 282882 121512 282888
rect 121458 282296 121514 282305
rect 121458 282231 121514 282240
rect 121472 281586 121500 282231
rect 121460 281580 121512 281586
rect 121460 281522 121512 281528
rect 121550 280936 121606 280945
rect 121550 280871 121606 280880
rect 121460 280288 121512 280294
rect 121458 280256 121460 280265
rect 121512 280256 121514 280265
rect 121564 280226 121592 280871
rect 121458 280191 121514 280200
rect 121552 280220 121604 280226
rect 121552 280162 121604 280168
rect 121550 279576 121606 279585
rect 121550 279511 121606 279520
rect 121458 278896 121514 278905
rect 121458 278831 121460 278840
rect 121512 278831 121514 278840
rect 121460 278802 121512 278808
rect 121564 278798 121592 279511
rect 121552 278792 121604 278798
rect 121552 278734 121604 278740
rect 121550 278216 121606 278225
rect 121550 278151 121606 278160
rect 121458 277536 121514 277545
rect 121458 277471 121460 277480
rect 121512 277471 121514 277480
rect 121460 277442 121512 277448
rect 121564 277438 121592 278151
rect 120828 277366 120948 277394
rect 121552 277432 121604 277438
rect 121552 277374 121604 277380
rect 120724 249552 120776 249558
rect 120724 249494 120776 249500
rect 120828 235754 120856 277366
rect 121460 277364 121512 277370
rect 121460 277306 121512 277312
rect 121472 276865 121500 277306
rect 121458 276856 121514 276865
rect 121458 276791 121514 276800
rect 121458 276176 121514 276185
rect 121458 276111 121514 276120
rect 121472 276078 121500 276111
rect 121460 276072 121512 276078
rect 121460 276014 121512 276020
rect 121656 275505 121684 309810
rect 122116 302190 122144 362238
rect 122104 302184 122156 302190
rect 122104 302126 122156 302132
rect 121734 290456 121790 290465
rect 121734 290391 121790 290400
rect 121748 289882 121776 290391
rect 121736 289876 121788 289882
rect 121736 289818 121788 289824
rect 122286 289096 122342 289105
rect 122286 289031 122342 289040
rect 121734 288416 121790 288425
rect 121734 288351 121790 288360
rect 121748 287094 121776 288351
rect 121736 287088 121788 287094
rect 121736 287030 121788 287036
rect 122300 286346 122328 289031
rect 122288 286340 122340 286346
rect 122288 286282 122340 286288
rect 121736 285660 121788 285666
rect 121736 285602 121788 285608
rect 121748 284345 121776 285602
rect 121734 284336 121790 284345
rect 121734 284271 121790 284280
rect 121734 281616 121790 281625
rect 121734 281551 121790 281560
rect 121748 279478 121776 281551
rect 121736 279472 121788 279478
rect 121736 279414 121788 279420
rect 121642 275496 121698 275505
rect 121642 275431 121698 275440
rect 121460 274644 121512 274650
rect 121460 274586 121512 274592
rect 121472 274145 121500 274586
rect 121458 274136 121514 274145
rect 121458 274071 121514 274080
rect 121656 273970 121684 275431
rect 121644 273964 121696 273970
rect 121644 273906 121696 273912
rect 121458 273456 121514 273465
rect 121458 273391 121514 273400
rect 121472 273290 121500 273391
rect 121460 273284 121512 273290
rect 121460 273226 121512 273232
rect 121552 273216 121604 273222
rect 121552 273158 121604 273164
rect 121564 272785 121592 273158
rect 121550 272776 121606 272785
rect 121550 272711 121606 272720
rect 122102 272096 122158 272105
rect 122102 272031 122158 272040
rect 121458 271416 121514 271425
rect 121458 271351 121514 271360
rect 121472 270570 121500 271351
rect 121460 270564 121512 270570
rect 121460 270506 121512 270512
rect 121642 270056 121698 270065
rect 121642 269991 121698 270000
rect 121458 269376 121514 269385
rect 121458 269311 121514 269320
rect 121472 269142 121500 269311
rect 121460 269136 121512 269142
rect 121460 269078 121512 269084
rect 121552 269068 121604 269074
rect 121552 269010 121604 269016
rect 121564 268705 121592 269010
rect 121550 268696 121606 268705
rect 121550 268631 121606 268640
rect 121656 268394 121684 269991
rect 121644 268388 121696 268394
rect 121644 268330 121696 268336
rect 121458 268016 121514 268025
rect 121458 267951 121514 267960
rect 121472 267782 121500 267951
rect 121460 267776 121512 267782
rect 121460 267718 121512 267724
rect 121550 267336 121606 267345
rect 121550 267271 121606 267280
rect 121458 266656 121514 266665
rect 121458 266591 121514 266600
rect 121472 266490 121500 266591
rect 121460 266484 121512 266490
rect 121460 266426 121512 266432
rect 121564 266422 121592 267271
rect 121552 266416 121604 266422
rect 121552 266358 121604 266364
rect 121550 265976 121606 265985
rect 121550 265911 121606 265920
rect 121458 265296 121514 265305
rect 121458 265231 121514 265240
rect 121472 265062 121500 265231
rect 121460 265056 121512 265062
rect 121460 264998 121512 265004
rect 121564 264994 121592 265911
rect 121552 264988 121604 264994
rect 121552 264930 121604 264936
rect 121460 264920 121512 264926
rect 121460 264862 121512 264868
rect 121472 264625 121500 264862
rect 121458 264616 121514 264625
rect 121458 264551 121514 264560
rect 121550 263936 121606 263945
rect 121550 263871 121606 263880
rect 121564 263634 121592 263871
rect 121552 263628 121604 263634
rect 121552 263570 121604 263576
rect 121460 263560 121512 263566
rect 121460 263502 121512 263508
rect 121472 263265 121500 263502
rect 121458 263256 121514 263265
rect 121458 263191 121514 263200
rect 121458 262576 121514 262585
rect 121458 262511 121514 262520
rect 121472 262274 121500 262511
rect 121460 262268 121512 262274
rect 121460 262210 121512 262216
rect 121550 261896 121606 261905
rect 121550 261831 121606 261840
rect 121564 260914 121592 261831
rect 121552 260908 121604 260914
rect 121552 260850 121604 260856
rect 121460 260840 121512 260846
rect 121460 260782 121512 260788
rect 121472 260545 121500 260782
rect 121458 260536 121514 260545
rect 121458 260471 121514 260480
rect 121458 259856 121514 259865
rect 121458 259791 121514 259800
rect 121472 259486 121500 259791
rect 121460 259480 121512 259486
rect 121460 259422 121512 259428
rect 121552 259412 121604 259418
rect 121552 259354 121604 259360
rect 121564 258505 121592 259354
rect 121642 259176 121698 259185
rect 121642 259111 121698 259120
rect 121550 258496 121606 258505
rect 121550 258431 121606 258440
rect 121656 258126 121684 259111
rect 121644 258120 121696 258126
rect 121644 258062 121696 258068
rect 121460 258052 121512 258058
rect 121460 257994 121512 258000
rect 121472 257145 121500 257994
rect 121550 257816 121606 257825
rect 121550 257751 121606 257760
rect 121458 257136 121514 257145
rect 121458 257071 121514 257080
rect 121564 256766 121592 257751
rect 121552 256760 121604 256766
rect 121552 256702 121604 256708
rect 121460 256692 121512 256698
rect 121460 256634 121512 256640
rect 121472 256465 121500 256634
rect 121552 256624 121604 256630
rect 121552 256566 121604 256572
rect 121458 256456 121514 256465
rect 121458 256391 121514 256400
rect 120908 256012 120960 256018
rect 120908 255954 120960 255960
rect 120920 238678 120948 255954
rect 121564 255785 121592 256566
rect 121550 255776 121606 255785
rect 121550 255711 121606 255720
rect 121550 255096 121606 255105
rect 121550 255031 121606 255040
rect 121458 254416 121514 254425
rect 121458 254351 121514 254360
rect 121472 254046 121500 254351
rect 121460 254040 121512 254046
rect 121460 253982 121512 253988
rect 121564 253978 121592 255031
rect 121552 253972 121604 253978
rect 121552 253914 121604 253920
rect 121550 253736 121606 253745
rect 121550 253671 121606 253680
rect 121458 253056 121514 253065
rect 121458 252991 121514 253000
rect 121472 252618 121500 252991
rect 121564 252686 121592 253671
rect 121552 252680 121604 252686
rect 121552 252622 121604 252628
rect 121460 252612 121512 252618
rect 121460 252554 121512 252560
rect 121458 251696 121514 251705
rect 121458 251631 121514 251640
rect 121472 251258 121500 251631
rect 121460 251252 121512 251258
rect 121460 251194 121512 251200
rect 121550 250336 121606 250345
rect 121550 250271 121606 250280
rect 121564 249830 121592 250271
rect 121552 249824 121604 249830
rect 121552 249766 121604 249772
rect 121460 249756 121512 249762
rect 121460 249698 121512 249704
rect 121472 249665 121500 249698
rect 121458 249656 121514 249665
rect 121458 249591 121514 249600
rect 121460 249552 121512 249558
rect 121460 249494 121512 249500
rect 121472 248402 121500 249494
rect 121550 248976 121606 248985
rect 121550 248911 121606 248920
rect 121564 248470 121592 248911
rect 121552 248464 121604 248470
rect 121552 248406 121604 248412
rect 121460 248396 121512 248402
rect 121460 248338 121512 248344
rect 121644 248396 121696 248402
rect 121644 248338 121696 248344
rect 121458 248296 121514 248305
rect 121458 248231 121514 248240
rect 121472 247110 121500 248231
rect 121656 247625 121684 248338
rect 121736 248328 121788 248334
rect 121736 248270 121788 248276
rect 121642 247616 121698 247625
rect 121642 247551 121698 247560
rect 121460 247104 121512 247110
rect 121460 247046 121512 247052
rect 121550 246936 121606 246945
rect 121550 246871 121606 246880
rect 121458 246256 121514 246265
rect 121458 246191 121514 246200
rect 121472 245682 121500 246191
rect 121564 245750 121592 246871
rect 121552 245744 121604 245750
rect 121552 245686 121604 245692
rect 121460 245676 121512 245682
rect 121460 245618 121512 245624
rect 121642 245576 121698 245585
rect 121642 245511 121698 245520
rect 121460 244248 121512 244254
rect 121460 244190 121512 244196
rect 121550 244216 121606 244225
rect 121472 243545 121500 244190
rect 121550 244151 121606 244160
rect 121458 243536 121514 243545
rect 121458 243471 121514 243480
rect 121564 242962 121592 244151
rect 121656 243574 121684 245511
rect 121748 244905 121776 248270
rect 121734 244896 121790 244905
rect 121734 244831 121790 244840
rect 121644 243568 121696 243574
rect 121644 243510 121696 243516
rect 121552 242956 121604 242962
rect 121552 242898 121604 242904
rect 121460 242888 121512 242894
rect 121458 242856 121460 242865
rect 121512 242856 121514 242865
rect 121458 242791 121514 242800
rect 121552 242820 121604 242826
rect 121552 242762 121604 242768
rect 121564 242185 121592 242762
rect 121550 242176 121606 242185
rect 121550 242111 121606 242120
rect 121460 241528 121512 241534
rect 121460 241470 121512 241476
rect 121472 240825 121500 241470
rect 121458 240816 121514 240825
rect 121458 240751 121514 240760
rect 121552 240780 121604 240786
rect 121552 240722 121604 240728
rect 121458 240136 121514 240145
rect 121458 240071 121514 240080
rect 121472 239766 121500 240071
rect 121460 239760 121512 239766
rect 121460 239702 121512 239708
rect 121564 238754 121592 240722
rect 121472 238726 121592 238754
rect 120908 238672 120960 238678
rect 120908 238614 120960 238620
rect 121472 238542 121500 238726
rect 121460 238536 121512 238542
rect 121460 238478 121512 238484
rect 120816 235748 120868 235754
rect 120816 235690 120868 235696
rect 120080 225616 120132 225622
rect 120080 225558 120132 225564
rect 115940 199504 115992 199510
rect 115940 199446 115992 199452
rect 119988 186380 120040 186386
rect 119988 186322 120040 186328
rect 114468 183592 114520 183598
rect 114468 183534 114520 183540
rect 112168 179444 112220 179450
rect 112168 179386 112220 179392
rect 112180 177041 112208 179386
rect 114480 177721 114508 183534
rect 116952 182300 117004 182306
rect 116952 182242 117004 182248
rect 115848 180940 115900 180946
rect 115848 180882 115900 180888
rect 115860 177721 115888 180882
rect 116964 177721 116992 182242
rect 120000 177721 120028 186322
rect 122116 181626 122144 272031
rect 122746 261216 122802 261225
rect 122852 261202 122880 380938
rect 123496 361554 123524 702714
rect 124864 630692 124916 630698
rect 124864 630634 124916 630640
rect 124220 385416 124272 385422
rect 124220 385358 124272 385364
rect 123484 361548 123536 361554
rect 123484 361490 123536 361496
rect 122932 358896 122984 358902
rect 122932 358838 122984 358844
rect 122802 261174 122880 261202
rect 122746 261151 122802 261160
rect 122944 241233 122972 358838
rect 123024 345160 123076 345166
rect 123024 345102 123076 345108
rect 123036 251054 123064 345102
rect 123116 305856 123168 305862
rect 123116 305798 123168 305804
rect 123128 263566 123156 305798
rect 124232 304298 124260 385358
rect 124876 339425 124904 630634
rect 126244 484424 126296 484430
rect 126244 484366 126296 484372
rect 125600 385280 125652 385286
rect 125600 385222 125652 385228
rect 124956 341556 125008 341562
rect 124956 341498 125008 341504
rect 124862 339416 124918 339425
rect 124862 339351 124918 339360
rect 124968 331226 124996 341498
rect 124312 331220 124364 331226
rect 124312 331162 124364 331168
rect 124956 331220 125008 331226
rect 124956 331162 125008 331168
rect 124220 304292 124272 304298
rect 124220 304234 124272 304240
rect 124220 302184 124272 302190
rect 124220 302126 124272 302132
rect 123116 263560 123168 263566
rect 123116 263502 123168 263508
rect 123024 251048 123076 251054
rect 123024 250990 123076 250996
rect 122930 241224 122986 241233
rect 122930 241159 122986 241168
rect 124232 238950 124260 302126
rect 124324 289814 124352 331162
rect 124404 316872 124456 316878
rect 124404 316814 124456 316820
rect 124416 312526 124444 316814
rect 124404 312520 124456 312526
rect 124404 312462 124456 312468
rect 124864 312520 124916 312526
rect 124864 312462 124916 312468
rect 124312 289808 124364 289814
rect 124312 289750 124364 289756
rect 124876 274650 124904 312462
rect 125048 294296 125100 294302
rect 125048 294238 125100 294244
rect 124864 274644 124916 274650
rect 124864 274586 124916 274592
rect 124956 272536 125008 272542
rect 124956 272478 125008 272484
rect 124864 239760 124916 239766
rect 124864 239702 124916 239708
rect 124220 238944 124272 238950
rect 124220 238886 124272 238892
rect 124876 195362 124904 239702
rect 124968 235686 124996 272478
rect 125060 265674 125088 294238
rect 125612 292534 125640 385222
rect 126256 339386 126284 484366
rect 130384 430636 130436 430642
rect 130384 430578 130436 430584
rect 128544 385212 128596 385218
rect 128544 385154 128596 385160
rect 128360 383988 128412 383994
rect 128360 383930 128412 383936
rect 127072 357468 127124 357474
rect 127072 357410 127124 357416
rect 125692 339380 125744 339386
rect 125692 339322 125744 339328
rect 126244 339380 126296 339386
rect 126244 339322 126296 339328
rect 125600 292528 125652 292534
rect 125600 292470 125652 292476
rect 125048 265668 125100 265674
rect 125048 265610 125100 265616
rect 125704 264926 125732 339322
rect 126980 336048 127032 336054
rect 126980 335990 127032 335996
rect 125876 297424 125928 297430
rect 125876 297366 125928 297372
rect 125782 293448 125838 293457
rect 125782 293383 125838 293392
rect 125796 285666 125824 293383
rect 125784 285660 125836 285666
rect 125784 285602 125836 285608
rect 125888 273222 125916 297366
rect 125876 273216 125928 273222
rect 125876 273158 125928 273164
rect 125692 264920 125744 264926
rect 125692 264862 125744 264868
rect 126992 256630 127020 335990
rect 127084 287026 127112 357410
rect 127164 298852 127216 298858
rect 127164 298794 127216 298800
rect 127072 287020 127124 287026
rect 127072 286962 127124 286968
rect 126980 256624 127032 256630
rect 126980 256566 127032 256572
rect 127176 238882 127204 298794
rect 127164 238876 127216 238882
rect 127164 238818 127216 238824
rect 124956 235680 125008 235686
rect 124956 235622 125008 235628
rect 128372 234530 128400 383930
rect 128452 376780 128504 376786
rect 128452 376722 128504 376728
rect 128464 242826 128492 376722
rect 128556 284306 128584 385154
rect 129740 351960 129792 351966
rect 129740 351902 129792 351908
rect 129004 317416 129056 317422
rect 129004 317358 129056 317364
rect 128544 284300 128596 284306
rect 128544 284242 128596 284248
rect 129016 258058 129044 317358
rect 129004 258052 129056 258058
rect 129004 257994 129056 258000
rect 128452 242820 128504 242826
rect 128452 242762 128504 242768
rect 129752 238746 129780 351902
rect 130396 338094 130424 430578
rect 136652 395350 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 700398 154160 703520
rect 154120 700392 154172 700398
rect 154120 700334 154172 700340
rect 155224 700392 155276 700398
rect 155224 700334 155276 700340
rect 142804 643136 142856 643142
rect 142804 643078 142856 643084
rect 141424 524476 141476 524482
rect 141424 524418 141476 524424
rect 136640 395344 136692 395350
rect 136640 395286 136692 395292
rect 135260 393984 135312 393990
rect 135260 393926 135312 393932
rect 135272 393378 135300 393926
rect 135260 393372 135312 393378
rect 135260 393314 135312 393320
rect 132500 386504 132552 386510
rect 132500 386446 132552 386452
rect 131212 380248 131264 380254
rect 131212 380190 131264 380196
rect 129832 338088 129884 338094
rect 129832 338030 129884 338036
rect 130384 338088 130436 338094
rect 130384 338030 130436 338036
rect 129844 256698 129872 338030
rect 131120 334756 131172 334762
rect 131120 334698 131172 334704
rect 129924 313948 129976 313954
rect 129924 313890 129976 313896
rect 129936 277370 129964 313890
rect 129924 277364 129976 277370
rect 129924 277306 129976 277312
rect 129936 276690 129964 277306
rect 129924 276684 129976 276690
rect 129924 276626 129976 276632
rect 129832 256692 129884 256698
rect 129832 256634 129884 256640
rect 131132 239018 131160 334698
rect 131224 317422 131252 380190
rect 131212 317416 131264 317422
rect 131212 317358 131264 317364
rect 132512 259418 132540 386446
rect 132592 383920 132644 383926
rect 132592 383862 132644 383868
rect 132604 269074 132632 383862
rect 133972 382424 134024 382430
rect 133972 382366 134024 382372
rect 133880 334688 133932 334694
rect 133880 334630 133932 334636
rect 132684 300144 132736 300150
rect 132684 300086 132736 300092
rect 132592 269068 132644 269074
rect 132592 269010 132644 269016
rect 132500 259412 132552 259418
rect 132500 259354 132552 259360
rect 132696 242894 132724 300086
rect 132684 242888 132736 242894
rect 132684 242830 132736 242836
rect 131120 239012 131172 239018
rect 131120 238954 131172 238960
rect 129740 238740 129792 238746
rect 129740 238682 129792 238688
rect 133892 235958 133920 334630
rect 133984 288386 134012 382366
rect 135168 349240 135220 349246
rect 135168 349182 135220 349188
rect 135180 348430 135208 349182
rect 135168 348424 135220 348430
rect 135168 348366 135220 348372
rect 134064 316804 134116 316810
rect 134064 316746 134116 316752
rect 133972 288380 134024 288386
rect 133972 288322 134024 288328
rect 134076 244254 134104 316746
rect 135168 288380 135220 288386
rect 135168 288322 135220 288328
rect 135180 287706 135208 288322
rect 135168 287700 135220 287706
rect 135168 287642 135220 287648
rect 134064 244248 134116 244254
rect 134064 244190 134116 244196
rect 135272 240786 135300 393314
rect 137100 388476 137152 388482
rect 137100 388418 137152 388424
rect 137112 387938 137140 388418
rect 136824 387932 136876 387938
rect 136824 387874 136876 387880
rect 137100 387932 137152 387938
rect 137100 387874 137152 387880
rect 136640 381064 136692 381070
rect 136640 381006 136692 381012
rect 135260 240780 135312 240786
rect 135260 240722 135312 240728
rect 133880 235952 133932 235958
rect 133880 235894 133932 235900
rect 135168 235952 135220 235958
rect 135168 235894 135220 235900
rect 135180 235278 135208 235894
rect 135168 235272 135220 235278
rect 135168 235214 135220 235220
rect 136652 234598 136680 381006
rect 136730 351928 136786 351937
rect 136730 351863 136786 351872
rect 136744 238610 136772 351863
rect 136836 286414 136864 387874
rect 140780 378208 140832 378214
rect 140780 378150 140832 378156
rect 139400 353320 139452 353326
rect 139400 353262 139452 353268
rect 136824 286408 136876 286414
rect 136824 286350 136876 286356
rect 139412 273222 139440 353262
rect 140792 293185 140820 378150
rect 141436 328438 141464 524418
rect 142160 364404 142212 364410
rect 142160 364346 142212 364352
rect 140872 328432 140924 328438
rect 140872 328374 140924 328380
rect 141424 328432 141476 328438
rect 141424 328374 141476 328380
rect 140778 293176 140834 293185
rect 140778 293111 140834 293120
rect 139400 273216 139452 273222
rect 139400 273158 139452 273164
rect 139412 272542 139440 273158
rect 139400 272536 139452 272542
rect 139400 272478 139452 272484
rect 140884 249762 140912 328374
rect 141424 295724 141476 295730
rect 141424 295666 141476 295672
rect 140872 249756 140924 249762
rect 140872 249698 140924 249704
rect 136732 238604 136784 238610
rect 136732 238546 136784 238552
rect 136640 234592 136692 234598
rect 136640 234534 136692 234540
rect 128360 234524 128412 234530
rect 128360 234466 128412 234472
rect 128372 233918 128400 234466
rect 128360 233912 128412 233918
rect 128360 233854 128412 233860
rect 133144 231192 133196 231198
rect 133144 231134 133196 231140
rect 133156 199578 133184 231134
rect 133144 199572 133196 199578
rect 133144 199514 133196 199520
rect 124864 195356 124916 195362
rect 124864 195298 124916 195304
rect 141436 188562 141464 295666
rect 142172 260846 142200 364346
rect 142816 351937 142844 643078
rect 146944 590708 146996 590714
rect 146944 590650 146996 590656
rect 142802 351928 142858 351937
rect 142802 351863 142858 351872
rect 146956 350606 146984 590650
rect 148324 563100 148376 563106
rect 148324 563042 148376 563048
rect 148336 389842 148364 563042
rect 148324 389836 148376 389842
rect 148324 389778 148376 389784
rect 155236 388482 155264 700334
rect 170324 700330 170352 703520
rect 202800 703186 202828 703520
rect 201500 703180 201552 703186
rect 201500 703122 201552 703128
rect 202788 703180 202840 703186
rect 202788 703122 202840 703128
rect 170312 700324 170364 700330
rect 170312 700266 170364 700272
rect 201512 391270 201540 703122
rect 218992 700398 219020 703520
rect 218980 700392 219032 700398
rect 218980 700334 219032 700340
rect 235184 700330 235212 703520
rect 220084 700324 220136 700330
rect 220084 700266 220136 700272
rect 235172 700324 235224 700330
rect 235172 700266 235224 700272
rect 220096 403646 220124 700266
rect 267660 697610 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 220084 403640 220136 403646
rect 220084 403582 220136 403588
rect 266372 393990 266400 697546
rect 282932 694822 282960 702406
rect 282920 694816 282972 694822
rect 282920 694758 282972 694764
rect 266360 393984 266412 393990
rect 266360 393926 266412 393932
rect 299492 392630 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703118 332548 703520
rect 332508 703112 332560 703118
rect 332508 703054 332560 703060
rect 348804 700330 348832 703520
rect 364996 703050 365024 703520
rect 364984 703044 365036 703050
rect 364984 702986 365036 702992
rect 341524 700324 341576 700330
rect 341524 700266 341576 700272
rect 348792 700324 348844 700330
rect 348792 700266 348844 700272
rect 299480 392624 299532 392630
rect 299480 392566 299532 392572
rect 201500 391264 201552 391270
rect 201500 391206 201552 391212
rect 166264 390584 166316 390590
rect 166264 390526 166316 390532
rect 155224 388476 155276 388482
rect 155224 388418 155276 388424
rect 147680 386572 147732 386578
rect 147680 386514 147732 386520
rect 143540 350600 143592 350606
rect 143540 350542 143592 350548
rect 146944 350600 146996 350606
rect 146944 350542 146996 350548
rect 142804 293276 142856 293282
rect 142804 293218 142856 293224
rect 142160 260840 142212 260846
rect 142160 260782 142212 260788
rect 142816 194002 142844 293218
rect 143448 260840 143500 260846
rect 143448 260782 143500 260788
rect 143460 260166 143488 260782
rect 143448 260160 143500 260166
rect 143448 260102 143500 260108
rect 143552 237386 143580 350542
rect 146944 315308 146996 315314
rect 146944 315250 146996 315256
rect 144184 298444 144236 298450
rect 144184 298386 144236 298392
rect 144092 276684 144144 276690
rect 144092 276626 144144 276632
rect 144104 269822 144132 276626
rect 144092 269816 144144 269822
rect 144092 269758 144144 269764
rect 143540 237380 143592 237386
rect 143540 237322 143592 237328
rect 142804 193996 142856 194002
rect 142804 193938 142856 193944
rect 144196 189854 144224 298386
rect 146956 192710 146984 315250
rect 147692 248402 147720 386514
rect 160744 385144 160796 385150
rect 160744 385086 160796 385092
rect 152464 326392 152516 326398
rect 152464 326334 152516 326340
rect 151084 302932 151136 302938
rect 151084 302874 151136 302880
rect 148324 278860 148376 278866
rect 148324 278802 148376 278808
rect 147680 248396 147732 248402
rect 147680 248338 147732 248344
rect 146944 192704 146996 192710
rect 146944 192646 146996 192652
rect 148336 191350 148364 278802
rect 148324 191344 148376 191350
rect 148324 191286 148376 191292
rect 144184 189848 144236 189854
rect 144184 189790 144236 189796
rect 141424 188556 141476 188562
rect 141424 188498 141476 188504
rect 129648 187808 129700 187814
rect 129648 187750 129700 187756
rect 128268 183660 128320 183666
rect 128268 183602 128320 183608
rect 122104 181620 122156 181626
rect 122104 181562 122156 181568
rect 120908 181008 120960 181014
rect 120908 180950 120960 180956
rect 120920 177721 120948 180950
rect 125416 179512 125468 179518
rect 125416 179454 125468 179460
rect 123300 178152 123352 178158
rect 123300 178094 123352 178100
rect 114466 177712 114522 177721
rect 114466 177647 114522 177656
rect 115846 177712 115902 177721
rect 115846 177647 115902 177656
rect 116950 177712 117006 177721
rect 116950 177647 117006 177656
rect 119986 177712 120042 177721
rect 119986 177647 120042 177656
rect 120906 177712 120962 177721
rect 120906 177647 120962 177656
rect 112166 177032 112222 177041
rect 112166 176967 112222 176976
rect 123312 176769 123340 178094
rect 125428 177041 125456 179454
rect 125414 177032 125470 177041
rect 125414 176967 125470 176976
rect 125876 176792 125928 176798
rect 123298 176760 123354 176769
rect 123298 176695 123354 176704
rect 125874 176760 125876 176769
rect 128280 176769 128308 183602
rect 129660 177721 129688 187750
rect 151096 185978 151124 302874
rect 152476 192778 152504 326334
rect 155224 319524 155276 319530
rect 155224 319466 155276 319472
rect 152464 192772 152516 192778
rect 152464 192714 152516 192720
rect 151084 185972 151136 185978
rect 151084 185914 151136 185920
rect 155236 183054 155264 319466
rect 159364 307148 159416 307154
rect 159364 307090 159416 307096
rect 155224 183048 155276 183054
rect 159376 183025 159404 307090
rect 155224 182990 155276 182996
rect 159362 183016 159418 183025
rect 159362 182951 159418 182960
rect 130752 180872 130804 180878
rect 130752 180814 130804 180820
rect 130764 177721 130792 180814
rect 160756 180266 160784 385086
rect 162122 379264 162178 379273
rect 162122 379199 162178 379208
rect 160744 180260 160796 180266
rect 160744 180202 160796 180208
rect 133144 178288 133196 178294
rect 133144 178230 133196 178236
rect 129646 177712 129702 177721
rect 129646 177647 129702 177656
rect 130750 177712 130806 177721
rect 130750 177647 130806 177656
rect 133156 176769 133184 178230
rect 148232 178220 148284 178226
rect 148232 178162 148284 178168
rect 134432 177064 134484 177070
rect 134432 177006 134484 177012
rect 134444 176769 134472 177006
rect 136088 176860 136140 176866
rect 136088 176802 136140 176808
rect 136100 176769 136128 176802
rect 148244 176769 148272 178162
rect 162136 177313 162164 379199
rect 166276 180334 166304 390526
rect 232504 389292 232556 389298
rect 232504 389234 232556 389240
rect 169024 387864 169076 387870
rect 169024 387806 169076 387812
rect 166354 302832 166410 302841
rect 166354 302767 166410 302776
rect 166264 180328 166316 180334
rect 166264 180270 166316 180276
rect 166368 180033 166396 302767
rect 166540 183660 166592 183666
rect 166540 183602 166592 183608
rect 166448 180940 166500 180946
rect 166448 180882 166500 180888
rect 166354 180024 166410 180033
rect 166354 179959 166410 179968
rect 164884 178288 164936 178294
rect 164884 178230 164936 178236
rect 162122 177304 162178 177313
rect 162122 177239 162178 177248
rect 125928 176760 125930 176769
rect 125874 176695 125930 176704
rect 128266 176760 128322 176769
rect 128266 176695 128322 176704
rect 133142 176760 133198 176769
rect 133142 176695 133198 176704
rect 134430 176760 134486 176769
rect 134430 176695 134486 176704
rect 136086 176760 136142 176769
rect 136086 176695 136142 176704
rect 148230 176760 148286 176769
rect 148230 176695 148286 176704
rect 132040 176316 132092 176322
rect 132040 176258 132092 176264
rect 118424 176180 118476 176186
rect 118424 176122 118476 176128
rect 111064 175976 111116 175982
rect 111064 175918 111116 175924
rect 118436 175409 118464 176122
rect 121920 176112 121972 176118
rect 121920 176054 121972 176060
rect 121932 175409 121960 176054
rect 127072 175976 127124 175982
rect 127072 175918 127124 175924
rect 127084 175545 127112 175918
rect 132052 175545 132080 176258
rect 158904 176248 158956 176254
rect 158904 176190 158956 176196
rect 158916 175545 158944 176190
rect 127070 175536 127126 175545
rect 127070 175471 127126 175480
rect 132038 175536 132094 175545
rect 132038 175471 132094 175480
rect 158902 175536 158958 175545
rect 158902 175471 158958 175480
rect 100758 175400 100814 175409
rect 100758 175335 100814 175344
rect 118422 175400 118478 175409
rect 118422 175335 118478 175344
rect 121918 175400 121974 175409
rect 121918 175335 121974 175344
rect 164896 175166 164924 178230
rect 166356 178152 166408 178158
rect 166356 178094 166408 178100
rect 165436 177064 165488 177070
rect 165436 177006 165488 177012
rect 165448 175234 165476 177006
rect 165528 176316 165580 176322
rect 165528 176258 165580 176264
rect 165436 175228 165488 175234
rect 165436 175170 165488 175176
rect 164884 175160 164936 175166
rect 164884 175102 164936 175108
rect 165540 173874 165568 176258
rect 166264 176180 166316 176186
rect 166264 176122 166316 176128
rect 165528 173868 165580 173874
rect 165528 173810 165580 173816
rect 166276 167006 166304 176122
rect 166368 169726 166396 178094
rect 166356 169720 166408 169726
rect 166356 169662 166408 169668
rect 166264 167000 166316 167006
rect 166264 166942 166316 166948
rect 166460 165578 166488 180882
rect 166552 172514 166580 183602
rect 167644 182232 167696 182238
rect 167644 182174 167696 182180
rect 166540 172508 166592 172514
rect 166540 172450 166592 172456
rect 166448 165572 166500 165578
rect 166448 165514 166500 165520
rect 167656 162858 167684 182174
rect 167736 181008 167788 181014
rect 167736 180950 167788 180956
rect 167748 168366 167776 180950
rect 167920 179512 167972 179518
rect 167920 179454 167972 179460
rect 167826 171592 167882 171601
rect 167826 171527 167882 171536
rect 167736 168360 167788 168366
rect 167736 168302 167788 168308
rect 167644 162852 167696 162858
rect 167644 162794 167696 162800
rect 167840 160750 167868 171527
rect 167932 169658 167960 179454
rect 167920 169652 167972 169658
rect 167920 169594 167972 169600
rect 167828 160744 167880 160750
rect 167828 160686 167880 160692
rect 167644 147688 167696 147694
rect 167644 147630 167696 147636
rect 166264 136672 166316 136678
rect 166264 136614 166316 136620
rect 66166 129296 66222 129305
rect 66166 129231 66222 129240
rect 65154 126304 65210 126313
rect 65154 126239 65210 126248
rect 65168 125662 65196 126239
rect 65156 125656 65208 125662
rect 65156 125598 65208 125604
rect 65522 125216 65578 125225
rect 65522 125151 65578 125160
rect 65536 124234 65564 125151
rect 65524 124228 65576 124234
rect 65524 124170 65576 124176
rect 66074 123584 66130 123593
rect 66074 123519 66130 123528
rect 66088 122874 66116 123519
rect 66076 122868 66128 122874
rect 66076 122810 66128 122816
rect 66074 102368 66130 102377
rect 66074 102303 66130 102312
rect 66088 81433 66116 102303
rect 66180 94897 66208 129231
rect 67454 128072 67510 128081
rect 67454 128007 67510 128016
rect 67362 122632 67418 122641
rect 67362 122567 67418 122576
rect 66166 94888 66222 94897
rect 66166 94823 66222 94832
rect 67376 91050 67404 122567
rect 67468 93809 67496 128007
rect 67546 120864 67602 120873
rect 67546 120799 67602 120808
rect 67454 93800 67510 93809
rect 67454 93735 67510 93744
rect 67364 91044 67416 91050
rect 67364 90986 67416 90992
rect 67560 84182 67588 120799
rect 67638 100736 67694 100745
rect 67638 100671 67694 100680
rect 67652 86970 67680 100671
rect 164884 98048 164936 98054
rect 164884 97990 164936 97996
rect 129370 94752 129426 94761
rect 129370 94687 129426 94696
rect 151726 94752 151782 94761
rect 151726 94687 151782 94696
rect 122840 94512 122892 94518
rect 122840 94454 122892 94460
rect 85670 93664 85726 93673
rect 85670 93599 85726 93608
rect 115478 93664 115534 93673
rect 115478 93599 115534 93608
rect 120630 93664 120686 93673
rect 120630 93599 120686 93608
rect 85684 93226 85712 93599
rect 115492 93294 115520 93599
rect 120644 93362 120672 93599
rect 120632 93356 120684 93362
rect 120632 93298 120684 93304
rect 115480 93288 115532 93294
rect 103426 93256 103482 93265
rect 85672 93220 85724 93226
rect 103426 93191 103482 93200
rect 110326 93256 110382 93265
rect 110326 93191 110382 93200
rect 113822 93256 113878 93265
rect 115480 93230 115532 93236
rect 113822 93191 113878 93200
rect 85672 93162 85724 93168
rect 74816 92472 74868 92478
rect 74814 92440 74816 92449
rect 74868 92440 74870 92449
rect 74814 92375 74870 92384
rect 88982 92440 89038 92449
rect 88982 92375 88984 92384
rect 89036 92375 89038 92384
rect 95054 92440 95110 92449
rect 95054 92375 95110 92384
rect 102046 92440 102102 92449
rect 102046 92375 102102 92384
rect 88984 92346 89036 92352
rect 95068 92342 95096 92375
rect 95056 92336 95108 92342
rect 95056 92278 95108 92284
rect 99194 91352 99250 91361
rect 99194 91287 99250 91296
rect 101862 91352 101918 91361
rect 101862 91287 101918 91296
rect 85486 91216 85542 91225
rect 85486 91151 85542 91160
rect 86866 91216 86922 91225
rect 86866 91151 86922 91160
rect 88062 91216 88118 91225
rect 88062 91151 88118 91160
rect 90730 91216 90786 91225
rect 90730 91151 90786 91160
rect 92386 91216 92442 91225
rect 92386 91151 92442 91160
rect 93766 91216 93822 91225
rect 93766 91151 93822 91160
rect 95146 91216 95202 91225
rect 95146 91151 95202 91160
rect 96526 91216 96582 91225
rect 96526 91151 96582 91160
rect 97078 91216 97134 91225
rect 97078 91151 97134 91160
rect 97906 91216 97962 91225
rect 97906 91151 97962 91160
rect 67640 86964 67692 86970
rect 67640 86906 67692 86912
rect 67548 84176 67600 84182
rect 67548 84118 67600 84124
rect 66074 81424 66130 81433
rect 66074 81359 66130 81368
rect 85500 77246 85528 91151
rect 86880 79898 86908 91151
rect 88076 86873 88104 91151
rect 90744 88262 90772 91151
rect 90732 88256 90784 88262
rect 90732 88198 90784 88204
rect 88062 86864 88118 86873
rect 88062 86799 88118 86808
rect 92400 81394 92428 91151
rect 92388 81388 92440 81394
rect 92388 81330 92440 81336
rect 86868 79892 86920 79898
rect 86868 79834 86920 79840
rect 93780 78538 93808 91151
rect 95160 79966 95188 91151
rect 96540 84046 96568 91151
rect 97092 86902 97120 91151
rect 97080 86896 97132 86902
rect 97080 86838 97132 86844
rect 96528 84040 96580 84046
rect 96528 83982 96580 83988
rect 95148 79960 95200 79966
rect 95148 79902 95200 79908
rect 97920 78674 97948 91151
rect 99208 82686 99236 91287
rect 99286 91216 99342 91225
rect 99286 91151 99342 91160
rect 100206 91216 100262 91225
rect 100206 91151 100262 91160
rect 100666 91216 100722 91225
rect 100666 91151 100722 91160
rect 99196 82680 99248 82686
rect 99196 82622 99248 82628
rect 99300 80073 99328 91151
rect 100220 88194 100248 91151
rect 100208 88188 100260 88194
rect 100208 88130 100260 88136
rect 100680 81258 100708 91151
rect 100668 81252 100720 81258
rect 100668 81194 100720 81200
rect 99286 80064 99342 80073
rect 99286 79999 99342 80008
rect 97908 78668 97960 78674
rect 97908 78610 97960 78616
rect 93768 78532 93820 78538
rect 93768 78474 93820 78480
rect 101876 78470 101904 91287
rect 101954 91216 102010 91225
rect 101954 91151 102010 91160
rect 101968 82618 101996 91151
rect 102060 91118 102088 92375
rect 102966 91216 103022 91225
rect 102966 91151 103022 91160
rect 102048 91112 102100 91118
rect 102048 91054 102100 91060
rect 102980 85542 103008 91151
rect 102968 85536 103020 85542
rect 102968 85478 103020 85484
rect 103440 84153 103468 93191
rect 105542 92440 105598 92449
rect 105542 92375 105598 92384
rect 106646 92440 106702 92449
rect 106646 92375 106702 92384
rect 105556 92274 105584 92375
rect 105544 92268 105596 92274
rect 105544 92210 105596 92216
rect 106094 91760 106150 91769
rect 106094 91695 106150 91704
rect 104806 91352 104862 91361
rect 104806 91287 104862 91296
rect 104714 91216 104770 91225
rect 104714 91151 104770 91160
rect 103426 84144 103482 84153
rect 103426 84079 103482 84088
rect 101956 82612 102008 82618
rect 101956 82554 102008 82560
rect 104728 81190 104756 91151
rect 104716 81184 104768 81190
rect 104716 81126 104768 81132
rect 101864 78464 101916 78470
rect 101864 78406 101916 78412
rect 85488 77240 85540 77246
rect 85488 77182 85540 77188
rect 92480 76560 92532 76566
rect 92480 76502 92532 76508
rect 69020 75200 69072 75206
rect 69020 75142 69072 75148
rect 67640 72480 67692 72486
rect 67640 72422 67692 72428
rect 64788 17400 64840 17406
rect 64788 17342 64840 17348
rect 60752 16546 60872 16574
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 60844 480 60872 16546
rect 62028 4820 62080 4826
rect 62028 4762 62080 4768
rect 62040 480 62068 4762
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 65524 6248 65576 6254
rect 65524 6190 65576 6196
rect 65536 480 65564 6190
rect 66720 2168 66772 2174
rect 66720 2110 66772 2116
rect 66732 480 66760 2110
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67652 354 67680 72422
rect 69032 6914 69060 75142
rect 71780 73840 71832 73846
rect 71780 73782 71832 73788
rect 70400 31068 70452 31074
rect 70400 31010 70452 31016
rect 69112 22840 69164 22846
rect 69112 22782 69164 22788
rect 69124 16574 69152 22782
rect 70412 16574 70440 31010
rect 71792 16574 71820 73782
rect 84200 72548 84252 72554
rect 84200 72490 84252 72496
rect 75920 69692 75972 69698
rect 75920 69634 75972 69640
rect 73160 46300 73212 46306
rect 73160 46242 73212 46248
rect 73172 16574 73200 46242
rect 74540 17264 74592 17270
rect 74540 17206 74592 17212
rect 74552 16574 74580 17206
rect 69124 16546 69888 16574
rect 70412 16546 71544 16574
rect 71792 16546 72648 16574
rect 73172 16546 73384 16574
rect 74552 16546 75040 16574
rect 69032 6886 69152 6914
rect 69124 480 69152 6886
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 16546
rect 71516 480 71544 16546
rect 72620 480 72648 16546
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75012 480 75040 16546
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 69634
rect 78680 68400 78732 68406
rect 78680 68342 78732 68348
rect 77300 32496 77352 32502
rect 77300 32438 77352 32444
rect 77312 6914 77340 32438
rect 77390 19952 77446 19961
rect 77390 19887 77446 19896
rect 77404 16574 77432 19887
rect 78692 16574 78720 68342
rect 82820 66972 82872 66978
rect 82820 66914 82872 66920
rect 81440 50448 81492 50454
rect 81440 50390 81492 50396
rect 81452 16574 81480 50390
rect 82832 16574 82860 66914
rect 77404 16546 78168 16574
rect 78692 16546 79272 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 77312 6886 77432 6914
rect 77404 480 77432 6886
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 79244 354 79272 16546
rect 80888 11756 80940 11762
rect 80888 11698 80940 11704
rect 80900 480 80928 11698
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 72490
rect 85580 65612 85632 65618
rect 85580 65554 85632 65560
rect 85592 3534 85620 65554
rect 89720 64184 89772 64190
rect 89720 64126 89772 64132
rect 88340 43512 88392 43518
rect 88340 43454 88392 43460
rect 85672 35216 85724 35222
rect 85672 35158 85724 35164
rect 85580 3528 85632 3534
rect 85580 3470 85632 3476
rect 85684 480 85712 35158
rect 86960 25628 87012 25634
rect 86960 25570 87012 25576
rect 86972 16574 87000 25570
rect 88352 16574 88380 43454
rect 89732 16574 89760 64126
rect 91100 19984 91152 19990
rect 91100 19926 91152 19932
rect 91112 16574 91140 19926
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 86500 3528 86552 3534
rect 86500 3470 86552 3476
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86512 354 86540 3470
rect 86838 354 86950 480
rect 86512 326 86950 354
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 76502
rect 104820 75886 104848 91287
rect 106108 89729 106136 91695
rect 106660 90914 106688 92375
rect 108210 91352 108266 91361
rect 108210 91287 108266 91296
rect 109590 91352 109646 91361
rect 109590 91287 109646 91296
rect 107198 91216 107254 91225
rect 107198 91151 107254 91160
rect 106648 90908 106700 90914
rect 106648 90850 106700 90856
rect 106094 89720 106150 89729
rect 106094 89655 106150 89664
rect 107212 88330 107240 91151
rect 107200 88324 107252 88330
rect 107200 88266 107252 88272
rect 108224 85474 108252 91287
rect 108486 91216 108542 91225
rect 108486 91151 108542 91160
rect 108500 86834 108528 91151
rect 108488 86828 108540 86834
rect 108488 86770 108540 86776
rect 108212 85468 108264 85474
rect 108212 85410 108264 85416
rect 109604 85406 109632 91287
rect 110142 91216 110198 91225
rect 110142 91151 110198 91160
rect 109592 85400 109644 85406
rect 109592 85342 109644 85348
rect 110156 82822 110184 91151
rect 110340 90846 110368 93191
rect 110694 91216 110750 91225
rect 110694 91151 110750 91160
rect 111706 91216 111762 91225
rect 111706 91151 111762 91160
rect 112534 91216 112590 91225
rect 112534 91151 112590 91160
rect 110328 90840 110380 90846
rect 110328 90782 110380 90788
rect 110708 88233 110736 91151
rect 110694 88224 110750 88233
rect 110694 88159 110750 88168
rect 111720 83978 111748 91151
rect 112548 85270 112576 91151
rect 113836 89622 113864 93191
rect 116766 92440 116822 92449
rect 116766 92375 116822 92384
rect 116780 92206 116808 92375
rect 122852 92342 122880 94454
rect 129384 93906 129412 94687
rect 151740 93974 151768 94687
rect 162860 94580 162912 94586
rect 162860 94522 162912 94528
rect 151728 93968 151780 93974
rect 151728 93910 151780 93916
rect 129372 93900 129424 93906
rect 129372 93842 129424 93848
rect 135718 93664 135774 93673
rect 135718 93599 135774 93608
rect 151726 93664 151782 93673
rect 151726 93599 151782 93608
rect 135732 93430 135760 93599
rect 151740 93498 151768 93599
rect 151728 93492 151780 93498
rect 151728 93434 151780 93440
rect 135720 93424 135772 93430
rect 135720 93366 135772 93372
rect 128174 93256 128230 93265
rect 128174 93191 128230 93200
rect 126612 93152 126664 93158
rect 126612 93094 126664 93100
rect 124034 92440 124090 92449
rect 124034 92375 124090 92384
rect 122840 92336 122892 92342
rect 122840 92278 122892 92284
rect 116768 92200 116820 92206
rect 116768 92142 116820 92148
rect 115570 91760 115626 91769
rect 115570 91695 115626 91704
rect 114466 91216 114522 91225
rect 114466 91151 114522 91160
rect 113824 89616 113876 89622
rect 113824 89558 113876 89564
rect 112536 85264 112588 85270
rect 112536 85206 112588 85212
rect 111708 83972 111760 83978
rect 111708 83914 111760 83920
rect 110144 82816 110196 82822
rect 110144 82758 110196 82764
rect 114480 77110 114508 91151
rect 115584 89690 115612 91695
rect 122838 91488 122894 91497
rect 122838 91423 122894 91432
rect 118238 91352 118294 91361
rect 118238 91287 118294 91296
rect 119894 91352 119950 91361
rect 119894 91287 119950 91296
rect 122654 91352 122710 91361
rect 122654 91287 122710 91296
rect 115846 91216 115902 91225
rect 115846 91151 115902 91160
rect 117134 91216 117190 91225
rect 117134 91151 117190 91160
rect 115572 89684 115624 89690
rect 115572 89626 115624 89632
rect 115860 84114 115888 91151
rect 117148 86766 117176 91151
rect 118252 88126 118280 91287
rect 118606 91216 118662 91225
rect 118606 91151 118662 91160
rect 118240 88120 118292 88126
rect 118240 88062 118292 88068
rect 117136 86760 117188 86766
rect 117136 86702 117188 86708
rect 115848 84108 115900 84114
rect 115848 84050 115900 84056
rect 118620 79830 118648 91151
rect 118700 91112 118752 91118
rect 118700 91054 118752 91060
rect 118712 89554 118740 91054
rect 118700 89548 118752 89554
rect 118700 89490 118752 89496
rect 119908 84017 119936 91287
rect 119986 91216 120042 91225
rect 119986 91151 120042 91160
rect 121366 91216 121422 91225
rect 121366 91151 121422 91160
rect 119894 84008 119950 84017
rect 119894 83943 119950 83952
rect 120000 80034 120028 91151
rect 119988 80028 120040 80034
rect 119988 79970 120040 79976
rect 118608 79824 118660 79830
rect 118608 79766 118660 79772
rect 121380 77178 121408 91151
rect 122668 82550 122696 91287
rect 122746 91216 122802 91225
rect 122746 91151 122802 91160
rect 122656 82544 122708 82550
rect 122656 82486 122708 82492
rect 122760 78606 122788 91151
rect 122852 85338 122880 91423
rect 124048 90778 124076 92375
rect 126624 92274 126652 93094
rect 126702 92440 126758 92449
rect 126702 92375 126758 92384
rect 126716 92274 126744 92375
rect 126612 92268 126664 92274
rect 126612 92210 126664 92216
rect 126704 92268 126756 92274
rect 126704 92210 126756 92216
rect 128188 92138 128216 93191
rect 134430 92440 134486 92449
rect 134430 92375 134486 92384
rect 153014 92440 153070 92449
rect 153014 92375 153070 92384
rect 134444 92342 134472 92375
rect 134432 92336 134484 92342
rect 134432 92278 134484 92284
rect 128176 92132 128228 92138
rect 128176 92074 128228 92080
rect 126702 92032 126758 92041
rect 126702 91967 126758 91976
rect 125414 91624 125470 91633
rect 125414 91559 125470 91568
rect 124126 91216 124182 91225
rect 124126 91151 124182 91160
rect 124036 90772 124088 90778
rect 124036 90714 124088 90720
rect 122840 85332 122892 85338
rect 122840 85274 122892 85280
rect 124140 82754 124168 91151
rect 125428 89418 125456 91559
rect 125506 91216 125562 91225
rect 125506 91151 125562 91160
rect 125416 89412 125468 89418
rect 125416 89354 125468 89360
rect 124128 82748 124180 82754
rect 124128 82690 124180 82696
rect 125520 81326 125548 91151
rect 126716 86698 126744 91967
rect 126886 91624 126942 91633
rect 126886 91559 126942 91568
rect 126900 89486 126928 91559
rect 131026 91216 131082 91225
rect 131026 91151 131082 91160
rect 132406 91216 132462 91225
rect 132406 91151 132462 91160
rect 133234 91216 133290 91225
rect 133234 91151 133290 91160
rect 151726 91216 151782 91225
rect 151726 91151 151782 91160
rect 126888 89480 126940 89486
rect 126888 89422 126940 89428
rect 126704 86692 126756 86698
rect 126704 86634 126756 86640
rect 125508 81320 125560 81326
rect 125508 81262 125560 81268
rect 131040 81122 131068 91151
rect 132420 88058 132448 91151
rect 132408 88052 132460 88058
rect 132408 87994 132460 88000
rect 133248 85202 133276 91151
rect 151740 90710 151768 91151
rect 151728 90704 151780 90710
rect 151728 90646 151780 90652
rect 153028 89350 153056 92375
rect 162872 89729 162900 94522
rect 164896 93226 164924 97990
rect 166276 93294 166304 136614
rect 166356 120148 166408 120154
rect 166356 120090 166408 120096
rect 166264 93288 166316 93294
rect 166264 93230 166316 93236
rect 164884 93220 164936 93226
rect 164884 93162 164936 93168
rect 162858 89720 162914 89729
rect 162858 89655 162914 89664
rect 153016 89344 153068 89350
rect 153016 89286 153068 89292
rect 166368 86766 166396 120090
rect 166448 110492 166500 110498
rect 166448 110434 166500 110440
rect 166460 88194 166488 110434
rect 166540 98116 166592 98122
rect 166540 98058 166592 98064
rect 166448 88188 166500 88194
rect 166448 88130 166500 88136
rect 166356 86760 166408 86766
rect 166356 86702 166408 86708
rect 133236 85196 133288 85202
rect 133236 85138 133288 85144
rect 131028 81116 131080 81122
rect 131028 81058 131080 81064
rect 166552 79898 166580 98058
rect 167656 93430 167684 147630
rect 167736 143608 167788 143614
rect 167736 143550 167788 143556
rect 167748 93906 167776 143550
rect 169036 115326 169064 387806
rect 195244 383784 195296 383790
rect 195244 383726 195296 383732
rect 173164 380180 173216 380186
rect 173164 380122 173216 380128
rect 169116 186516 169168 186522
rect 169116 186458 169168 186464
rect 169128 157350 169156 186458
rect 171784 186448 171836 186454
rect 171784 186390 171836 186396
rect 169300 183592 169352 183598
rect 169300 183534 169352 183540
rect 169208 176996 169260 177002
rect 169208 176938 169260 176944
rect 169220 158710 169248 176938
rect 169312 165510 169340 183534
rect 170588 182300 170640 182306
rect 170588 182242 170640 182248
rect 170496 179444 170548 179450
rect 170496 179386 170548 179392
rect 170404 178084 170456 178090
rect 170404 178026 170456 178032
rect 169300 165504 169352 165510
rect 169300 165446 169352 165452
rect 170416 162790 170444 178026
rect 170508 164218 170536 179386
rect 170600 166938 170628 182242
rect 171140 181620 171192 181626
rect 171140 181562 171192 181568
rect 170680 176112 170732 176118
rect 170680 176054 170732 176060
rect 170692 168298 170720 176054
rect 170680 168292 170732 168298
rect 170680 168234 170732 168240
rect 170588 166932 170640 166938
rect 170588 166874 170640 166880
rect 170496 164212 170548 164218
rect 170496 164154 170548 164160
rect 170404 162784 170456 162790
rect 170404 162726 170456 162732
rect 169208 158704 169260 158710
rect 169208 158646 169260 158652
rect 169116 157344 169168 157350
rect 169116 157286 169168 157292
rect 169208 124228 169260 124234
rect 169208 124170 169260 124176
rect 169116 122868 169168 122874
rect 169116 122810 169168 122816
rect 169024 115320 169076 115326
rect 169024 115262 169076 115268
rect 168288 111784 168340 111790
rect 168286 111752 168288 111761
rect 168340 111752 168342 111761
rect 168286 111687 168342 111696
rect 167828 110424 167880 110430
rect 167828 110366 167880 110372
rect 167840 110129 167868 110366
rect 167826 110120 167882 110129
rect 167826 110055 167882 110064
rect 169024 109064 169076 109070
rect 169024 109006 169076 109012
rect 168104 108996 168156 109002
rect 168104 108938 168156 108944
rect 168116 108769 168144 108938
rect 168102 108760 168158 108769
rect 168102 108695 168158 108704
rect 167828 106344 167880 106350
rect 167828 106286 167880 106292
rect 167736 93900 167788 93906
rect 167736 93842 167788 93848
rect 167644 93424 167696 93430
rect 167644 93366 167696 93372
rect 166540 79892 166592 79898
rect 166540 79834 166592 79840
rect 122748 78600 122800 78606
rect 122748 78542 122800 78548
rect 167840 78538 167868 106286
rect 167920 97300 167972 97306
rect 167920 97242 167972 97248
rect 167932 92410 167960 97242
rect 167920 92404 167972 92410
rect 167920 92346 167972 92352
rect 169036 84046 169064 109006
rect 169024 84040 169076 84046
rect 169024 83982 169076 83988
rect 169128 82550 169156 122810
rect 169220 90778 169248 124170
rect 170588 122936 170640 122942
rect 170588 122878 170640 122884
rect 170404 118856 170456 118862
rect 170404 118798 170456 118804
rect 169300 101448 169352 101454
rect 169300 101390 169352 101396
rect 169312 92206 169340 101390
rect 169300 92200 169352 92206
rect 169300 92142 169352 92148
rect 169208 90772 169260 90778
rect 169208 90714 169260 90720
rect 170416 85270 170444 118798
rect 170496 111852 170548 111858
rect 170496 111794 170548 111800
rect 170404 85264 170456 85270
rect 170404 85206 170456 85212
rect 169116 82544 169168 82550
rect 169116 82486 169168 82492
rect 170508 81258 170536 111794
rect 170600 93362 170628 122878
rect 170680 117360 170732 117366
rect 170680 117302 170732 117308
rect 170588 93356 170640 93362
rect 170588 93298 170640 93304
rect 170692 90846 170720 117302
rect 170680 90840 170732 90846
rect 170680 90782 170732 90788
rect 170496 81252 170548 81258
rect 170496 81194 170548 81200
rect 167828 78532 167880 78538
rect 167828 78474 167880 78480
rect 121368 77172 121420 77178
rect 121368 77114 121420 77120
rect 114468 77104 114520 77110
rect 114468 77046 114520 77052
rect 104808 75880 104860 75886
rect 104808 75822 104860 75828
rect 95240 75268 95292 75274
rect 95240 75210 95292 75216
rect 93860 62824 93912 62830
rect 93860 62766 93912 62772
rect 93872 6914 93900 62766
rect 93952 46232 94004 46238
rect 93952 46174 94004 46180
rect 93964 16574 93992 46174
rect 95252 16574 95280 75210
rect 122840 73976 122892 73982
rect 122840 73918 122892 73924
rect 99380 73908 99432 73914
rect 99380 73850 99432 73856
rect 98000 71120 98052 71126
rect 98000 71062 98052 71068
rect 96620 61464 96672 61470
rect 96620 61406 96672 61412
rect 96632 16574 96660 61406
rect 98012 16574 98040 71062
rect 99392 16574 99420 73850
rect 115940 72616 115992 72622
rect 115940 72558 115992 72564
rect 110420 69760 110472 69766
rect 110420 69702 110472 69708
rect 100760 58744 100812 58750
rect 100760 58686 100812 58692
rect 93964 16546 94728 16574
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 93872 6886 93992 6914
rect 93964 480 93992 6886
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 58686
rect 103520 57316 103572 57322
rect 103520 57258 103572 57264
rect 102140 24132 102192 24138
rect 102140 24074 102192 24080
rect 102152 16574 102180 24074
rect 103532 16574 103560 57258
rect 107660 55956 107712 55962
rect 107660 55898 107712 55904
rect 106280 49156 106332 49162
rect 106280 49098 106332 49104
rect 106292 16574 106320 49098
rect 107672 16574 107700 55898
rect 109040 35284 109092 35290
rect 109040 35226 109092 35232
rect 102152 16546 102272 16574
rect 103532 16546 104112 16574
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 102244 480 102272 16546
rect 103336 3528 103388 3534
rect 103336 3470 103388 3476
rect 103348 480 103376 3470
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105728 7608 105780 7614
rect 105728 7550 105780 7556
rect 105740 480 105768 7550
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109052 354 109080 35226
rect 110432 6914 110460 69702
rect 113180 68468 113232 68474
rect 113180 68410 113232 68416
rect 110512 54596 110564 54602
rect 110512 54538 110564 54544
rect 110524 16574 110552 54538
rect 111800 17332 111852 17338
rect 111800 17274 111852 17280
rect 111812 16574 111840 17274
rect 113192 16574 113220 68410
rect 114560 53100 114612 53106
rect 114560 53042 114612 53048
rect 114572 16574 114600 53042
rect 115952 16574 115980 72558
rect 121460 49088 121512 49094
rect 121460 49030 121512 49036
rect 118700 26988 118752 26994
rect 118700 26930 118752 26936
rect 118712 16574 118740 26930
rect 120080 25696 120132 25702
rect 120080 25638 120132 25644
rect 120092 16574 120120 25638
rect 121472 16574 121500 49030
rect 122852 16574 122880 73918
rect 124220 51808 124272 51814
rect 124220 51750 124272 51756
rect 124232 16574 124260 51750
rect 110524 16546 111656 16574
rect 111812 16546 112392 16574
rect 113192 16546 114048 16574
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 118712 16546 118832 16574
rect 120092 16546 120672 16574
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 124232 16546 124720 16574
rect 110432 6886 110552 6914
rect 110524 480 110552 6886
rect 111628 480 111656 16546
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114020 480 114048 16546
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 117596 4888 117648 4894
rect 117596 4830 117648 4836
rect 117608 480 117636 4830
rect 118804 480 118832 16546
rect 119896 9036 119948 9042
rect 119896 8978 119948 8984
rect 119908 480 119936 8978
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 122300 480 122328 16546
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124692 480 124720 16546
rect 168380 7676 168432 7682
rect 168380 7618 168432 7624
rect 125876 3596 125928 3602
rect 125876 3538 125928 3544
rect 125888 480 125916 3538
rect 168392 480 168420 7618
rect 171152 3602 171180 181562
rect 171796 155922 171824 186390
rect 171784 155916 171836 155922
rect 171784 155858 171836 155864
rect 171784 140820 171836 140826
rect 171784 140762 171836 140768
rect 171796 89418 171824 140762
rect 171876 131164 171928 131170
rect 171876 131106 171928 131112
rect 171784 89412 171836 89418
rect 171784 89354 171836 89360
rect 171888 81190 171916 131106
rect 171968 129804 172020 129810
rect 171968 129746 172020 129752
rect 171980 82618 172008 129746
rect 173176 104174 173204 380122
rect 186964 358828 187016 358834
rect 186964 358770 187016 358776
rect 180064 311160 180116 311166
rect 180064 311102 180116 311108
rect 178682 294128 178738 294137
rect 178682 294063 178738 294072
rect 177304 285728 177356 285734
rect 177304 285670 177356 285676
rect 177316 247722 177344 285670
rect 177304 247716 177356 247722
rect 177304 247658 177356 247664
rect 177304 187808 177356 187814
rect 177304 187750 177356 187756
rect 173256 187740 173308 187746
rect 173256 187682 173308 187688
rect 173268 160070 173296 187682
rect 177316 172446 177344 187750
rect 177304 172440 177356 172446
rect 177304 172382 177356 172388
rect 173256 160064 173308 160070
rect 173256 160006 173308 160012
rect 175924 153264 175976 153270
rect 175924 153206 175976 153212
rect 174544 146328 174596 146334
rect 174544 146270 174596 146276
rect 173256 142180 173308 142186
rect 173256 142122 173308 142128
rect 173164 104168 173216 104174
rect 173164 104110 173216 104116
rect 173164 100768 173216 100774
rect 173164 100710 173216 100716
rect 171968 82612 172020 82618
rect 171968 82554 172020 82560
rect 171876 81184 171928 81190
rect 171876 81126 171928 81132
rect 173176 77246 173204 100710
rect 173268 86698 173296 142122
rect 173348 132524 173400 132530
rect 173348 132466 173400 132472
rect 173360 90914 173388 132466
rect 173440 115252 173492 115258
rect 173440 115194 173492 115200
rect 173452 92138 173480 115194
rect 173440 92132 173492 92138
rect 173440 92074 173492 92080
rect 173348 90908 173400 90914
rect 173348 90850 173400 90856
rect 173256 86692 173308 86698
rect 173256 86634 173308 86640
rect 174556 85202 174584 146270
rect 174636 144968 174688 144974
rect 174636 144910 174688 144916
rect 174648 88058 174676 144910
rect 174728 117428 174780 117434
rect 174728 117370 174780 117376
rect 174636 88052 174688 88058
rect 174636 87994 174688 88000
rect 174544 85196 174596 85202
rect 174544 85138 174596 85144
rect 174740 83978 174768 117370
rect 175936 93498 175964 153206
rect 177304 151836 177356 151842
rect 177304 151778 177356 151784
rect 176016 128376 176068 128382
rect 176016 128318 176068 128324
rect 175924 93492 175976 93498
rect 175924 93434 175976 93440
rect 174728 83972 174780 83978
rect 174728 83914 174780 83920
rect 176028 78470 176056 128318
rect 176108 125656 176160 125662
rect 176108 125598 176160 125604
rect 176120 89486 176148 125598
rect 177316 90710 177344 151778
rect 177580 137284 177632 137290
rect 177580 137226 177632 137232
rect 177396 121508 177448 121514
rect 177396 121450 177448 121456
rect 177304 90704 177356 90710
rect 177304 90646 177356 90652
rect 176108 89480 176160 89486
rect 176108 89422 176160 89428
rect 177408 88126 177436 121450
rect 177488 110560 177540 110566
rect 177488 110502 177540 110508
rect 177396 88120 177448 88126
rect 177396 88062 177448 88068
rect 177500 82686 177528 110502
rect 177592 110430 177620 137226
rect 177580 110424 177632 110430
rect 177580 110366 177632 110372
rect 177580 106412 177632 106418
rect 177580 106354 177632 106360
rect 177488 82680 177540 82686
rect 177488 82622 177540 82628
rect 177592 81394 177620 106354
rect 178696 95169 178724 294063
rect 178868 153332 178920 153338
rect 178868 153274 178920 153280
rect 178776 135312 178828 135318
rect 178776 135254 178828 135260
rect 178682 95160 178738 95169
rect 178682 95095 178738 95104
rect 178684 91792 178736 91798
rect 178684 91734 178736 91740
rect 177580 81388 177632 81394
rect 177580 81330 177632 81336
rect 176016 78464 176068 78470
rect 176016 78406 176068 78412
rect 173164 77240 173216 77246
rect 173164 77182 173216 77188
rect 171140 3596 171192 3602
rect 171140 3538 171192 3544
rect 178696 3466 178724 91734
rect 178788 77110 178816 135254
rect 178880 93974 178908 153274
rect 178960 108316 179012 108322
rect 178960 108258 179012 108264
rect 178868 93968 178920 93974
rect 178868 93910 178920 93916
rect 178972 92313 179000 108258
rect 178958 92304 179014 92313
rect 178958 92239 179014 92248
rect 180076 77994 180104 311102
rect 184204 238128 184256 238134
rect 184204 238070 184256 238076
rect 180156 235272 180208 235278
rect 180156 235214 180208 235220
rect 180064 77988 180116 77994
rect 180064 77930 180116 77936
rect 178776 77104 178828 77110
rect 178776 77046 178828 77052
rect 180168 46918 180196 235214
rect 182824 180328 182876 180334
rect 182824 180270 182876 180276
rect 181444 178220 181496 178226
rect 181444 178162 181496 178168
rect 181456 150414 181484 178162
rect 181444 150408 181496 150414
rect 181444 150350 181496 150356
rect 180340 140072 180392 140078
rect 180340 140014 180392 140020
rect 180248 113212 180300 113218
rect 180248 113154 180300 113160
rect 180260 75886 180288 113154
rect 180352 109002 180380 140014
rect 181444 133952 181496 133958
rect 181444 133894 181496 133900
rect 180340 108996 180392 109002
rect 180340 108938 180392 108944
rect 181456 85406 181484 133894
rect 181536 116000 181588 116006
rect 181536 115942 181588 115948
rect 181548 86834 181576 115942
rect 181536 86828 181588 86834
rect 181536 86770 181588 86776
rect 181444 85400 181496 85406
rect 181444 85342 181496 85348
rect 180248 75880 180300 75886
rect 180248 75822 180300 75828
rect 180156 46912 180208 46918
rect 180156 46854 180208 46860
rect 182836 28354 182864 180270
rect 184216 177342 184244 238070
rect 184204 177336 184256 177342
rect 184204 177278 184256 177284
rect 185582 177304 185638 177313
rect 185582 177239 185638 177248
rect 184848 176928 184900 176934
rect 184848 176870 184900 176876
rect 184860 176050 184888 176870
rect 184204 176044 184256 176050
rect 184204 175986 184256 175992
rect 184848 176044 184900 176050
rect 184848 175986 184900 175992
rect 184216 157282 184244 175986
rect 184204 157276 184256 157282
rect 184204 157218 184256 157224
rect 184296 151904 184348 151910
rect 184296 151846 184348 151852
rect 184204 145036 184256 145042
rect 184204 144978 184256 144984
rect 182916 107704 182968 107710
rect 182916 107646 182968 107652
rect 182928 79966 182956 107646
rect 184216 81122 184244 144978
rect 184308 89350 184336 151846
rect 184296 89344 184348 89350
rect 184296 89286 184348 89292
rect 184204 81116 184256 81122
rect 184204 81058 184256 81064
rect 182916 79960 182968 79966
rect 182916 79902 182968 79908
rect 185596 60110 185624 177239
rect 185676 118788 185728 118794
rect 185676 118730 185728 118736
rect 185688 89622 185716 118730
rect 185676 89616 185728 89622
rect 185676 89558 185728 89564
rect 185584 60104 185636 60110
rect 185584 60046 185636 60052
rect 182824 28348 182876 28354
rect 182824 28290 182876 28296
rect 186976 10470 187004 358770
rect 191104 337544 191156 337550
rect 191104 337486 191156 337492
rect 188344 337476 188396 337482
rect 188344 337418 188396 337424
rect 187056 185972 187108 185978
rect 187056 185914 187108 185920
rect 187068 11898 187096 185914
rect 187148 124296 187200 124302
rect 187148 124238 187200 124244
rect 187160 85338 187188 124238
rect 188356 89010 188384 337418
rect 188436 189100 188488 189106
rect 188436 189042 188488 189048
rect 188448 161430 188476 189042
rect 189722 180024 189778 180033
rect 189722 179959 189778 179968
rect 188436 161424 188488 161430
rect 188436 161366 188488 161372
rect 188436 120216 188488 120222
rect 188436 120158 188488 120164
rect 188344 89004 188396 89010
rect 188344 88946 188396 88952
rect 188344 87644 188396 87650
rect 188344 87586 188396 87592
rect 187148 85332 187200 85338
rect 187148 85274 187200 85280
rect 187056 11892 187108 11898
rect 187056 11834 187108 11840
rect 186964 10464 187016 10470
rect 186964 10406 187016 10412
rect 188356 3534 188384 87586
rect 188448 84114 188476 120158
rect 188528 104916 188580 104922
rect 188528 104858 188580 104864
rect 188540 88262 188568 104858
rect 188528 88256 188580 88262
rect 188528 88198 188580 88204
rect 188436 84108 188488 84114
rect 188436 84050 188488 84056
rect 189736 21554 189764 179959
rect 189816 111920 189868 111926
rect 189816 111862 189868 111868
rect 189828 89554 189856 111862
rect 189816 89548 189868 89554
rect 189816 89490 189868 89496
rect 189724 21548 189776 21554
rect 189724 21490 189776 21496
rect 191116 18766 191144 337486
rect 192484 300960 192536 300966
rect 192484 300902 192536 300908
rect 192496 191282 192524 300902
rect 192484 191276 192536 191282
rect 192484 191218 192536 191224
rect 193864 183048 193916 183054
rect 191194 183016 191250 183025
rect 193864 182990 193916 182996
rect 191194 182951 191250 182960
rect 191104 18760 191156 18766
rect 191104 18702 191156 18708
rect 191208 11830 191236 182951
rect 192484 180260 192536 180266
rect 192484 180202 192536 180208
rect 192496 14618 192524 180202
rect 192576 103556 192628 103562
rect 192576 103498 192628 103504
rect 192588 90982 192616 103498
rect 192576 90976 192628 90982
rect 192576 90918 192628 90924
rect 193876 24206 193904 182990
rect 195256 29782 195284 383726
rect 215944 383716 215996 383722
rect 215944 383658 215996 383664
rect 209044 382696 209096 382702
rect 209044 382638 209096 382644
rect 196624 374060 196676 374066
rect 196624 374002 196676 374008
rect 195336 294160 195388 294166
rect 195336 294102 195388 294108
rect 195348 93673 195376 294102
rect 195520 109132 195572 109138
rect 195520 109074 195572 109080
rect 195426 106856 195482 106865
rect 195426 106791 195482 106800
rect 195334 93664 195390 93673
rect 195334 93599 195390 93608
rect 195244 29776 195296 29782
rect 195244 29718 195296 29724
rect 193864 24200 193916 24206
rect 193864 24142 193916 24148
rect 195440 16046 195468 106791
rect 195532 78674 195560 109074
rect 196636 83502 196664 374002
rect 202144 360324 202196 360330
rect 202144 360266 202196 360272
rect 198004 319456 198056 319462
rect 198004 319398 198056 319404
rect 196716 138032 196768 138038
rect 196716 137974 196768 137980
rect 196624 83496 196676 83502
rect 196624 83438 196676 83444
rect 196728 79830 196756 137974
rect 196716 79824 196768 79830
rect 196716 79766 196768 79772
rect 195520 78668 195572 78674
rect 195520 78610 195572 78616
rect 195428 16040 195480 16046
rect 195428 15982 195480 15988
rect 192484 14612 192536 14618
rect 192484 14554 192536 14560
rect 191196 11824 191248 11830
rect 191196 11766 191248 11772
rect 198016 7682 198044 319398
rect 199384 301028 199436 301034
rect 199384 300970 199436 300976
rect 199396 192642 199424 300970
rect 200764 192772 200816 192778
rect 200764 192714 200816 192720
rect 199384 192636 199436 192642
rect 199384 192578 199436 192584
rect 199476 189780 199528 189786
rect 199476 189722 199528 189728
rect 198096 176248 198148 176254
rect 198096 176190 198148 176196
rect 198108 149054 198136 176190
rect 198096 149048 198148 149054
rect 198096 148990 198148 148996
rect 198096 127016 198148 127022
rect 198096 126958 198148 126964
rect 198108 86902 198136 126958
rect 198188 116068 198240 116074
rect 198188 116010 198240 116016
rect 198096 86896 198148 86902
rect 198096 86838 198148 86844
rect 198200 82822 198228 116010
rect 199382 115152 199438 115161
rect 199382 115087 199438 115096
rect 198188 82816 198240 82822
rect 198188 82758 198240 82764
rect 198004 7676 198056 7682
rect 198004 7618 198056 7624
rect 199396 6322 199424 115087
rect 199488 96626 199516 189722
rect 199568 150476 199620 150482
rect 199568 150418 199620 150424
rect 199580 111790 199608 150418
rect 199568 111784 199620 111790
rect 199568 111726 199620 111732
rect 199568 102196 199620 102202
rect 199568 102138 199620 102144
rect 199476 96620 199528 96626
rect 199476 96562 199528 96568
rect 199580 93537 199608 102138
rect 199566 93528 199622 93537
rect 199566 93463 199622 93472
rect 200776 9110 200804 192714
rect 202156 86290 202184 360266
rect 206284 354748 206336 354754
rect 206284 354690 206336 354696
rect 204904 327752 204956 327758
rect 204904 327694 204956 327700
rect 202236 296948 202288 296954
rect 202236 296890 202288 296896
rect 202248 188630 202276 296890
rect 203524 295588 203576 295594
rect 203524 295530 203576 295536
rect 202236 188624 202288 188630
rect 202236 188566 202288 188572
rect 203536 187066 203564 295530
rect 203524 187060 203576 187066
rect 203524 187002 203576 187008
rect 202236 176724 202288 176730
rect 202236 176666 202288 176672
rect 202248 158642 202276 176666
rect 202236 158636 202288 158642
rect 202236 158578 202288 158584
rect 202236 142248 202288 142254
rect 202236 142190 202288 142196
rect 202248 92274 202276 142190
rect 202328 132592 202380 132598
rect 202328 132534 202380 132540
rect 202236 92268 202288 92274
rect 202236 92210 202288 92216
rect 202144 86284 202196 86290
rect 202144 86226 202196 86232
rect 202340 85474 202368 132534
rect 203616 131232 203668 131238
rect 203616 131174 203668 131180
rect 203524 115320 203576 115326
rect 203524 115262 203576 115268
rect 202328 85468 202380 85474
rect 202328 85410 202380 85416
rect 203536 13122 203564 115262
rect 203628 94586 203656 131174
rect 203708 102264 203760 102270
rect 203708 102206 203760 102212
rect 203616 94580 203668 94586
rect 203616 94522 203668 94528
rect 203720 91050 203748 102206
rect 203708 91044 203760 91050
rect 203708 90986 203760 90992
rect 203524 13116 203576 13122
rect 203524 13058 203576 13064
rect 200764 9104 200816 9110
rect 200764 9046 200816 9052
rect 199384 6316 199436 6322
rect 199384 6258 199436 6264
rect 188344 3528 188396 3534
rect 188344 3470 188396 3476
rect 204916 3466 204944 327694
rect 204996 318096 205048 318102
rect 204996 318038 205048 318044
rect 205008 24274 205036 318038
rect 206296 84862 206324 354690
rect 206376 347812 206428 347818
rect 206376 347754 206428 347760
rect 206284 84856 206336 84862
rect 206284 84798 206336 84804
rect 206388 82142 206416 347754
rect 207664 296880 207716 296886
rect 207664 296822 207716 296828
rect 207676 181626 207704 296822
rect 207664 181620 207716 181626
rect 207664 181562 207716 181568
rect 207664 139460 207716 139466
rect 207664 139402 207716 139408
rect 206560 103624 206612 103630
rect 206560 103566 206612 103572
rect 206468 100836 206520 100842
rect 206468 100778 206520 100784
rect 206480 84182 206508 100778
rect 206572 95062 206600 103566
rect 206560 95056 206612 95062
rect 206560 94998 206612 95004
rect 206468 84176 206520 84182
rect 206468 84118 206520 84124
rect 206376 82136 206428 82142
rect 206376 82078 206428 82084
rect 207676 77178 207704 139402
rect 207756 125724 207808 125730
rect 207756 125666 207808 125672
rect 207768 81326 207796 125666
rect 207756 81320 207808 81326
rect 207756 81262 207808 81268
rect 209056 80714 209084 382638
rect 211804 356108 211856 356114
rect 211804 356050 211856 356056
rect 210516 298376 210568 298382
rect 210516 298318 210568 298324
rect 209228 292868 209280 292874
rect 209228 292810 209280 292816
rect 209136 192704 209188 192710
rect 209136 192646 209188 192652
rect 209044 80708 209096 80714
rect 209044 80650 209096 80656
rect 207664 77172 207716 77178
rect 207664 77114 207716 77120
rect 204996 24268 205048 24274
rect 204996 24210 205048 24216
rect 209148 15978 209176 192646
rect 209240 188698 209268 292810
rect 210424 248464 210476 248470
rect 210424 248406 210476 248412
rect 209228 188692 209280 188698
rect 209228 188634 209280 188640
rect 209228 121576 209280 121582
rect 209228 121518 209280 121524
rect 209240 80034 209268 121518
rect 210436 95198 210464 248406
rect 210528 185609 210556 298318
rect 210514 185600 210570 185609
rect 210514 185535 210570 185544
rect 210608 146396 210660 146402
rect 210608 146338 210660 146344
rect 210516 140888 210568 140894
rect 210516 140830 210568 140836
rect 210424 95192 210476 95198
rect 210424 95134 210476 95140
rect 210528 82754 210556 140830
rect 210620 92342 210648 146338
rect 210608 92336 210660 92342
rect 210608 92278 210660 92284
rect 210516 82748 210568 82754
rect 210516 82690 210568 82696
rect 209228 80028 209280 80034
rect 209228 79970 209280 79976
rect 211816 78062 211844 356050
rect 213184 316736 213236 316742
rect 213184 316678 213236 316684
rect 211896 175976 211948 175982
rect 211896 175918 211948 175924
rect 211908 171086 211936 175918
rect 211896 171080 211948 171086
rect 211896 171022 211948 171028
rect 211896 114572 211948 114578
rect 211896 114514 211948 114520
rect 211908 88330 211936 114514
rect 211896 88324 211948 88330
rect 211896 88266 211948 88272
rect 211804 78056 211856 78062
rect 211804 77998 211856 78004
rect 209136 15972 209188 15978
rect 209136 15914 209188 15920
rect 213196 3602 213224 316678
rect 213276 299804 213328 299810
rect 213276 299746 213328 299752
rect 213288 189922 213316 299746
rect 214564 273284 214616 273290
rect 214564 273226 214616 273232
rect 213276 189916 213328 189922
rect 213276 189858 213328 189864
rect 214576 178838 214604 273226
rect 214656 227044 214708 227050
rect 214656 226986 214708 226992
rect 214668 184414 214696 226986
rect 214748 186380 214800 186386
rect 214748 186322 214800 186328
rect 214656 184408 214708 184414
rect 214656 184350 214708 184356
rect 214656 180872 214708 180878
rect 214656 180814 214708 180820
rect 214564 178832 214616 178838
rect 214564 178774 214616 178780
rect 213920 176860 213972 176866
rect 213920 176802 213972 176808
rect 213932 176225 213960 176802
rect 213918 176216 213974 176225
rect 213918 176151 213974 176160
rect 214564 176044 214616 176050
rect 214564 175986 214616 175992
rect 213920 175228 213972 175234
rect 213920 175170 213972 175176
rect 213932 175137 213960 175170
rect 214012 175160 214064 175166
rect 213918 175128 213974 175137
rect 214012 175102 214064 175108
rect 213918 175063 213974 175072
rect 214024 174729 214052 175102
rect 214010 174720 214066 174729
rect 214010 174655 214066 174664
rect 213920 173868 213972 173874
rect 213920 173810 213972 173816
rect 213932 173777 213960 173810
rect 213918 173768 213974 173777
rect 213918 173703 213974 173712
rect 214012 172508 214064 172514
rect 214012 172450 214064 172456
rect 213920 172440 213972 172446
rect 213918 172408 213920 172417
rect 213972 172408 213974 172417
rect 213918 172343 213974 172352
rect 214024 172009 214052 172450
rect 214010 172000 214066 172009
rect 214010 171935 214066 171944
rect 214576 171134 214604 175986
rect 214668 173369 214696 180814
rect 214654 173360 214710 173369
rect 214654 173295 214710 173304
rect 214576 171106 214696 171134
rect 214472 171080 214524 171086
rect 214472 171022 214524 171028
rect 214484 170921 214512 171022
rect 214470 170912 214526 170921
rect 214470 170847 214526 170856
rect 214012 169720 214064 169726
rect 213918 169688 213974 169697
rect 214012 169662 214064 169668
rect 213918 169623 213920 169632
rect 213972 169623 213974 169632
rect 213920 169594 213972 169600
rect 214024 169425 214052 169662
rect 214010 169416 214066 169425
rect 214010 169351 214066 169360
rect 214012 168360 214064 168366
rect 213918 168328 213974 168337
rect 214012 168302 214064 168308
rect 213918 168263 213920 168272
rect 213972 168263 213974 168272
rect 213920 168234 213972 168240
rect 214024 168065 214052 168302
rect 214010 168056 214066 168065
rect 214010 167991 214066 168000
rect 214012 167000 214064 167006
rect 214012 166942 214064 166948
rect 213920 166932 213972 166938
rect 213920 166874 213972 166880
rect 213932 166161 213960 166874
rect 214024 166705 214052 166942
rect 214010 166696 214066 166705
rect 214010 166631 214066 166640
rect 213918 166152 213974 166161
rect 213918 166087 213974 166096
rect 213920 165572 213972 165578
rect 213920 165514 213972 165520
rect 213932 165345 213960 165514
rect 214012 165504 214064 165510
rect 214012 165446 214064 165452
rect 213918 165336 213974 165345
rect 213918 165271 213974 165280
rect 214024 164801 214052 165446
rect 214010 164792 214066 164801
rect 214010 164727 214066 164736
rect 213920 164212 213972 164218
rect 213920 164154 213972 164160
rect 213932 163441 213960 164154
rect 213918 163432 213974 163441
rect 213918 163367 213974 163376
rect 213920 162852 213972 162858
rect 213920 162794 213972 162800
rect 213932 162625 213960 162794
rect 214012 162784 214064 162790
rect 214012 162726 214064 162732
rect 213918 162616 213974 162625
rect 213918 162551 213974 162560
rect 214024 162081 214052 162726
rect 214010 162072 214066 162081
rect 214010 162007 214066 162016
rect 213920 161424 213972 161430
rect 213920 161366 213972 161372
rect 213932 160857 213960 161366
rect 214668 161265 214696 171106
rect 214760 166977 214788 186322
rect 214932 176792 214984 176798
rect 214932 176734 214984 176740
rect 214944 170785 214972 176734
rect 214930 170776 214986 170785
rect 214930 170711 214986 170720
rect 214746 166968 214802 166977
rect 214746 166903 214802 166912
rect 214654 161256 214710 161265
rect 214654 161191 214710 161200
rect 213918 160848 213974 160857
rect 213918 160783 213974 160792
rect 214656 160744 214708 160750
rect 214656 160686 214708 160692
rect 213920 160064 213972 160070
rect 213920 160006 213972 160012
rect 213932 158817 213960 160006
rect 213918 158808 213974 158817
rect 213918 158743 213974 158752
rect 213920 158704 213972 158710
rect 213918 158672 213920 158681
rect 213972 158672 213974 158681
rect 213918 158607 213974 158616
rect 214012 158636 214064 158642
rect 214012 158578 214064 158584
rect 214024 158137 214052 158578
rect 214010 158128 214066 158137
rect 214010 158063 214066 158072
rect 214012 157344 214064 157350
rect 213918 157312 213974 157321
rect 214012 157286 214064 157292
rect 213918 157247 213920 157256
rect 213972 157247 213974 157256
rect 213920 157218 213972 157224
rect 214024 156913 214052 157286
rect 214010 156904 214066 156913
rect 214010 156839 214066 156848
rect 213918 155952 213974 155961
rect 213918 155887 213920 155896
rect 213972 155887 213974 155896
rect 213920 155858 213972 155864
rect 214010 153912 214066 153921
rect 214010 153847 214066 153856
rect 213918 153504 213974 153513
rect 213918 153439 213974 153448
rect 213932 153270 213960 153439
rect 214024 153338 214052 153847
rect 214012 153332 214064 153338
rect 214012 153274 214064 153280
rect 213920 153264 213972 153270
rect 213920 153206 213972 153212
rect 214010 152688 214066 152697
rect 214010 152623 214066 152632
rect 213918 152008 213974 152017
rect 213918 151943 213974 151952
rect 213932 151910 213960 151943
rect 213920 151904 213972 151910
rect 213920 151846 213972 151852
rect 214024 151842 214052 152623
rect 214562 151872 214618 151881
rect 214012 151836 214064 151842
rect 214562 151807 214618 151816
rect 214012 151778 214064 151784
rect 213918 150648 213974 150657
rect 213918 150583 213974 150592
rect 213932 150482 213960 150583
rect 213920 150476 213972 150482
rect 213920 150418 213972 150424
rect 214012 150408 214064 150414
rect 214012 150350 214064 150356
rect 214024 150113 214052 150350
rect 214010 150104 214066 150113
rect 214010 150039 214066 150048
rect 213920 149048 213972 149054
rect 213920 148990 213972 148996
rect 213932 148753 213960 148990
rect 213918 148744 213974 148753
rect 213918 148679 213974 148688
rect 213918 148064 213974 148073
rect 213918 147999 213974 148008
rect 213932 147694 213960 147999
rect 213920 147688 213972 147694
rect 213920 147630 213972 147636
rect 214010 146704 214066 146713
rect 214010 146639 214066 146648
rect 213918 146432 213974 146441
rect 214024 146402 214052 146639
rect 213918 146367 213974 146376
rect 214012 146396 214064 146402
rect 213932 146334 213960 146367
rect 214012 146338 214064 146344
rect 213920 146328 213972 146334
rect 213920 146270 213972 146276
rect 214010 145344 214066 145353
rect 214010 145279 214066 145288
rect 213920 145036 213972 145042
rect 213920 144978 213972 144984
rect 213932 144945 213960 144978
rect 214024 144974 214052 145279
rect 214012 144968 214064 144974
rect 213918 144936 213974 144945
rect 214012 144910 214064 144916
rect 213918 144871 213974 144880
rect 213918 143984 213974 143993
rect 213918 143919 213974 143928
rect 213932 143614 213960 143919
rect 213920 143608 213972 143614
rect 213920 143550 213972 143556
rect 214010 142760 214066 142769
rect 214010 142695 214066 142704
rect 213918 142352 213974 142361
rect 213918 142287 213974 142296
rect 213932 142254 213960 142287
rect 213920 142248 213972 142254
rect 213920 142190 213972 142196
rect 214024 142186 214052 142695
rect 214012 142180 214064 142186
rect 214012 142122 214064 142128
rect 213918 141400 213974 141409
rect 213918 141335 213974 141344
rect 213932 140826 213960 141335
rect 214010 140992 214066 141001
rect 214010 140927 214066 140936
rect 214024 140894 214052 140927
rect 214012 140888 214064 140894
rect 214012 140830 214064 140836
rect 213920 140820 213972 140826
rect 213920 140762 213972 140768
rect 214576 140078 214604 151807
rect 214668 149569 214696 160686
rect 214746 150784 214802 150793
rect 214746 150719 214802 150728
rect 214654 149560 214710 149569
rect 214654 149495 214710 149504
rect 214760 142154 214788 150719
rect 214838 143576 214894 143585
rect 214838 143511 214894 143520
rect 214668 142126 214788 142154
rect 214564 140072 214616 140078
rect 213274 140040 213330 140049
rect 214564 140014 214616 140020
rect 213274 139975 213330 139984
rect 213288 78606 213316 139975
rect 213918 139496 213974 139505
rect 213918 139431 213920 139440
rect 213972 139431 213974 139440
rect 213920 139402 213972 139408
rect 213918 138136 213974 138145
rect 213918 138071 213974 138080
rect 213932 138038 213960 138071
rect 213920 138032 213972 138038
rect 213920 137974 213972 137980
rect 214470 137456 214526 137465
rect 214668 137442 214696 142126
rect 214470 137391 214526 137400
rect 214576 137414 214696 137442
rect 213918 136776 213974 136785
rect 213918 136711 213974 136720
rect 213932 136678 213960 136711
rect 213920 136672 213972 136678
rect 213920 136614 213972 136620
rect 213918 135688 213974 135697
rect 213918 135623 213974 135632
rect 213932 135318 213960 135623
rect 213920 135312 213972 135318
rect 213920 135254 213972 135260
rect 213918 134056 213974 134065
rect 213918 133991 213974 134000
rect 213932 133958 213960 133991
rect 213920 133952 213972 133958
rect 213920 133894 213972 133900
rect 214010 132832 214066 132841
rect 214010 132767 214066 132776
rect 214024 132598 214052 132767
rect 214012 132592 214064 132598
rect 213918 132560 213974 132569
rect 214012 132534 214064 132540
rect 213918 132495 213920 132504
rect 213972 132495 213974 132504
rect 213920 132466 213972 132472
rect 214484 132494 214512 137391
rect 214576 137290 214604 137414
rect 214852 137306 214880 143511
rect 214564 137284 214616 137290
rect 214564 137226 214616 137232
rect 214668 137278 214880 137306
rect 214484 132466 214604 132494
rect 214010 131472 214066 131481
rect 214010 131407 214066 131416
rect 214024 131238 214052 131407
rect 214012 131232 214064 131238
rect 213918 131200 213974 131209
rect 214012 131174 214064 131180
rect 213918 131135 213920 131144
rect 213972 131135 213974 131144
rect 213920 131106 213972 131112
rect 213918 129840 213974 129849
rect 213918 129775 213920 129784
rect 213972 129775 213974 129784
rect 213920 129746 213972 129752
rect 213918 128888 213974 128897
rect 213918 128823 213974 128832
rect 213932 128382 213960 128823
rect 213920 128376 213972 128382
rect 213920 128318 213972 128324
rect 213918 127120 213974 127129
rect 213918 127055 213974 127064
rect 213932 127022 213960 127055
rect 213920 127016 213972 127022
rect 213920 126958 213972 126964
rect 214010 126168 214066 126177
rect 214010 126103 214066 126112
rect 213918 125760 213974 125769
rect 213918 125695 213920 125704
rect 213972 125695 213974 125704
rect 213920 125666 213972 125672
rect 214024 125662 214052 126103
rect 214012 125656 214064 125662
rect 214012 125598 214064 125604
rect 214010 124808 214066 124817
rect 214010 124743 214066 124752
rect 213918 124400 213974 124409
rect 213918 124335 213974 124344
rect 213932 124302 213960 124335
rect 213920 124296 213972 124302
rect 213920 124238 213972 124244
rect 214024 124234 214052 124743
rect 214012 124228 214064 124234
rect 214012 124170 214064 124176
rect 214010 123584 214066 123593
rect 214010 123519 214066 123528
rect 213918 123176 213974 123185
rect 213918 123111 213974 123120
rect 213932 122942 213960 123111
rect 213920 122936 213972 122942
rect 213920 122878 213972 122884
rect 214024 122874 214052 123519
rect 214012 122868 214064 122874
rect 214012 122810 214064 122816
rect 214010 122224 214066 122233
rect 214010 122159 214066 122168
rect 214024 121582 214052 122159
rect 214012 121576 214064 121582
rect 213918 121544 213974 121553
rect 214012 121518 214064 121524
rect 213918 121479 213920 121488
rect 213972 121479 213974 121488
rect 213920 121450 213972 121456
rect 214010 120864 214066 120873
rect 214010 120799 214066 120808
rect 213918 120456 213974 120465
rect 213918 120391 213974 120400
rect 213932 120222 213960 120391
rect 213920 120216 213972 120222
rect 213920 120158 213972 120164
rect 214024 120154 214052 120799
rect 214012 120148 214064 120154
rect 214012 120090 214064 120096
rect 213366 119640 213422 119649
rect 213366 119575 213422 119584
rect 213380 89690 213408 119575
rect 214010 119096 214066 119105
rect 214010 119031 214066 119040
rect 213918 118960 213974 118969
rect 213918 118895 213974 118904
rect 213932 118862 213960 118895
rect 213920 118856 213972 118862
rect 213920 118798 213972 118804
rect 214024 118794 214052 119031
rect 214012 118788 214064 118794
rect 214012 118730 214064 118736
rect 214010 117600 214066 117609
rect 214010 117535 214066 117544
rect 214024 117434 214052 117535
rect 214012 117428 214064 117434
rect 214012 117370 214064 117376
rect 213920 117360 213972 117366
rect 213918 117328 213920 117337
rect 213972 117328 213974 117337
rect 213918 117263 213974 117272
rect 214010 116240 214066 116249
rect 214010 116175 214066 116184
rect 214024 116074 214052 116175
rect 214012 116068 214064 116074
rect 214012 116010 214064 116016
rect 213920 116000 213972 116006
rect 213918 115968 213920 115977
rect 213972 115968 213974 115977
rect 213918 115903 213974 115912
rect 213918 115016 213974 115025
rect 213918 114951 213974 114960
rect 213932 114578 213960 114951
rect 213920 114572 213972 114578
rect 213920 114514 213972 114520
rect 213918 113656 213974 113665
rect 213918 113591 213974 113600
rect 213458 113248 213514 113257
rect 213932 113218 213960 113591
rect 213458 113183 213514 113192
rect 213920 113212 213972 113218
rect 213368 89684 213420 89690
rect 213368 89626 213420 89632
rect 213472 85542 213500 113183
rect 213920 113154 213972 113160
rect 214010 112296 214066 112305
rect 214010 112231 214066 112240
rect 214024 111926 214052 112231
rect 214012 111920 214064 111926
rect 213918 111888 213974 111897
rect 214012 111862 214064 111868
rect 213918 111823 213920 111832
rect 213972 111823 213974 111832
rect 213920 111794 213972 111800
rect 214010 110936 214066 110945
rect 214010 110871 214066 110880
rect 213920 110560 213972 110566
rect 213918 110528 213920 110537
rect 213972 110528 213974 110537
rect 214024 110498 214052 110871
rect 213918 110463 213974 110472
rect 214012 110492 214064 110498
rect 214012 110434 214064 110440
rect 214010 109712 214066 109721
rect 214010 109647 214066 109656
rect 213918 109304 213974 109313
rect 213918 109239 213974 109248
rect 213932 109070 213960 109239
rect 214024 109138 214052 109647
rect 214012 109132 214064 109138
rect 214012 109074 214064 109080
rect 213920 109064 213972 109070
rect 213920 109006 213972 109012
rect 213918 107944 213974 107953
rect 213918 107879 213974 107888
rect 213932 107710 213960 107879
rect 213920 107704 213972 107710
rect 213920 107646 213972 107652
rect 214010 106992 214066 107001
rect 214010 106927 214066 106936
rect 213918 106448 213974 106457
rect 213918 106383 213920 106392
rect 213972 106383 213974 106392
rect 213920 106354 213972 106360
rect 214024 106350 214052 106927
rect 214012 106344 214064 106350
rect 214012 106286 214064 106292
rect 213918 105768 213974 105777
rect 213918 105703 213974 105712
rect 213932 104922 213960 105703
rect 213920 104916 213972 104922
rect 213920 104858 213972 104864
rect 214010 104000 214066 104009
rect 214010 103935 214066 103944
rect 213918 103728 213974 103737
rect 213918 103663 213974 103672
rect 213932 103562 213960 103663
rect 214024 103630 214052 103935
rect 214012 103624 214064 103630
rect 214012 103566 214064 103572
rect 213920 103556 213972 103562
rect 214576 103514 214604 132466
rect 214668 115258 214696 137278
rect 214746 136096 214802 136105
rect 214746 136031 214802 136040
rect 214656 115252 214708 115258
rect 214656 115194 214708 115200
rect 214654 108352 214710 108361
rect 214760 108322 214788 136031
rect 215022 114608 215078 114617
rect 215022 114543 215078 114552
rect 214654 108287 214710 108296
rect 214748 108316 214800 108322
rect 213920 103498 213972 103504
rect 214484 103486 214604 103514
rect 214010 102504 214066 102513
rect 214010 102439 214066 102448
rect 213918 102368 213974 102377
rect 213918 102303 213974 102312
rect 213932 102270 213960 102303
rect 213920 102264 213972 102270
rect 213920 102206 213972 102212
rect 214024 102202 214052 102439
rect 214012 102196 214064 102202
rect 214012 102138 214064 102144
rect 214484 101454 214512 103486
rect 214472 101448 214524 101454
rect 214472 101390 214524 101396
rect 214010 101280 214066 101289
rect 214010 101215 214066 101224
rect 213918 101144 213974 101153
rect 213918 101079 213974 101088
rect 213932 100774 213960 101079
rect 214024 100842 214052 101215
rect 214012 100836 214064 100842
rect 214012 100778 214064 100784
rect 213920 100768 213972 100774
rect 213920 100710 213972 100716
rect 214102 99784 214158 99793
rect 214102 99719 214158 99728
rect 214010 98424 214066 98433
rect 214010 98359 214066 98368
rect 214024 98122 214052 98359
rect 214012 98116 214064 98122
rect 214012 98058 214064 98064
rect 213920 98048 213972 98054
rect 213918 98016 213920 98025
rect 213972 98016 213974 98025
rect 213918 97951 213974 97960
rect 214116 97306 214144 99719
rect 214104 97300 214156 97306
rect 214104 97242 214156 97248
rect 214562 96656 214618 96665
rect 214562 96591 214618 96600
rect 214576 86970 214604 96591
rect 214668 94518 214696 108287
rect 214748 108258 214800 108264
rect 215036 103514 215064 114543
rect 214852 103486 215064 103514
rect 214746 95840 214802 95849
rect 214746 95775 214802 95784
rect 214656 94512 214708 94518
rect 214656 94454 214708 94460
rect 214760 92478 214788 95775
rect 214852 93158 214880 103486
rect 214840 93152 214892 93158
rect 214840 93094 214892 93100
rect 214748 92472 214800 92478
rect 214748 92414 214800 92420
rect 214564 86964 214616 86970
rect 214564 86906 214616 86912
rect 213460 85536 213512 85542
rect 213460 85478 213512 85484
rect 213276 78600 213328 78606
rect 213276 78542 213328 78548
rect 213184 3596 213236 3602
rect 213184 3538 213236 3544
rect 215956 3534 215984 383658
rect 216036 345092 216088 345098
rect 216036 345034 216088 345040
rect 216048 7750 216076 345034
rect 217324 305652 217376 305658
rect 217324 305594 217376 305600
rect 216128 292800 216180 292806
rect 216128 292742 216180 292748
rect 216140 95130 216168 292742
rect 216220 104168 216272 104174
rect 216220 104110 216272 104116
rect 216128 95124 216180 95130
rect 216128 95066 216180 95072
rect 216232 13190 216260 104110
rect 216220 13184 216272 13190
rect 216220 13126 216272 13132
rect 216036 7744 216088 7750
rect 216036 7686 216088 7692
rect 217336 3670 217364 305594
rect 229744 303748 229796 303754
rect 229744 303690 229796 303696
rect 226984 303680 227036 303686
rect 226984 303622 227036 303628
rect 222844 302388 222896 302394
rect 222844 302330 222896 302336
rect 218704 294228 218756 294234
rect 218704 294170 218756 294176
rect 218716 192545 218744 294170
rect 220084 256760 220136 256766
rect 220084 256702 220136 256708
rect 218702 192536 218758 192545
rect 218702 192471 218758 192480
rect 220096 180266 220124 256702
rect 222856 183054 222884 302330
rect 224224 300892 224276 300898
rect 224224 300834 224276 300840
rect 222936 289944 222988 289950
rect 222936 289886 222988 289892
rect 222844 183048 222896 183054
rect 222844 182990 222896 182996
rect 222948 180334 222976 289886
rect 224236 183190 224264 300834
rect 224316 245744 224368 245750
rect 224316 245686 224368 245692
rect 224224 183184 224276 183190
rect 224224 183126 224276 183132
rect 222936 180328 222988 180334
rect 222936 180270 222988 180276
rect 220084 180260 220136 180266
rect 220084 180202 220136 180208
rect 224328 177410 224356 245686
rect 226996 183122 227024 303622
rect 227076 280288 227128 280294
rect 227076 280230 227128 280236
rect 226984 183116 227036 183122
rect 226984 183058 227036 183064
rect 227088 178906 227116 280230
rect 228364 224324 228416 224330
rect 228364 224266 228416 224272
rect 227076 178900 227128 178906
rect 227076 178842 227128 178848
rect 228376 177478 228404 224266
rect 229756 186969 229784 303690
rect 231124 292732 231176 292738
rect 231124 292674 231176 292680
rect 229742 186960 229798 186969
rect 229742 186895 229798 186904
rect 228364 177472 228416 177478
rect 231136 177449 231164 292674
rect 231216 245676 231268 245682
rect 231216 245618 231268 245624
rect 231228 181762 231256 245618
rect 231216 181756 231268 181762
rect 231216 181698 231268 181704
rect 228364 177414 228416 177420
rect 231122 177440 231178 177449
rect 224316 177404 224368 177410
rect 231122 177375 231178 177384
rect 224316 177346 224368 177352
rect 232516 177313 232544 389234
rect 313924 386436 313976 386442
rect 313924 386378 313976 386384
rect 309784 385076 309836 385082
rect 309784 385018 309836 385024
rect 280804 382628 280856 382634
rect 280804 382570 280856 382576
rect 271880 370524 271932 370530
rect 271880 370466 271932 370472
rect 269764 349172 269816 349178
rect 269764 349114 269816 349120
rect 269120 336184 269172 336190
rect 269120 336126 269172 336132
rect 246304 306468 246356 306474
rect 246304 306410 246356 306416
rect 244924 302456 244976 302462
rect 244924 302398 244976 302404
rect 232596 299736 232648 299742
rect 232596 299678 232648 299684
rect 232608 185978 232636 299678
rect 238024 299668 238076 299674
rect 238024 299610 238076 299616
rect 233884 269136 233936 269142
rect 233884 269078 233936 269084
rect 232596 185972 232648 185978
rect 232596 185914 232648 185920
rect 233896 177546 233924 269078
rect 233976 263628 234028 263634
rect 233976 263570 234028 263576
rect 233988 180402 234016 263570
rect 235264 259480 235316 259486
rect 235264 259422 235316 259428
rect 233976 180396 234028 180402
rect 233976 180338 234028 180344
rect 235276 178974 235304 259422
rect 236644 210520 236696 210526
rect 236644 210462 236696 210468
rect 235264 178968 235316 178974
rect 235264 178910 235316 178916
rect 233884 177540 233936 177546
rect 233884 177482 233936 177488
rect 232502 177304 232558 177313
rect 232502 177239 232558 177248
rect 236656 175982 236684 210462
rect 238036 181694 238064 299610
rect 240784 295452 240836 295458
rect 240784 295394 240836 295400
rect 238116 249824 238168 249830
rect 238116 249766 238168 249772
rect 238024 181688 238076 181694
rect 238024 181630 238076 181636
rect 238128 176254 238156 249766
rect 239404 202292 239456 202298
rect 239404 202234 239456 202240
rect 239416 180470 239444 202234
rect 239496 191344 239548 191350
rect 239496 191286 239548 191292
rect 239404 180464 239456 180470
rect 239404 180406 239456 180412
rect 238116 176248 238168 176254
rect 238116 176190 238168 176196
rect 239508 176186 239536 191286
rect 240796 178809 240824 295394
rect 240876 281580 240928 281586
rect 240876 281522 240928 281528
rect 240782 178800 240838 178809
rect 240782 178735 240838 178744
rect 240888 177585 240916 281522
rect 242164 221536 242216 221542
rect 242164 221478 242216 221484
rect 242176 178022 242204 221478
rect 242256 189848 242308 189854
rect 242256 189790 242308 189796
rect 242164 178016 242216 178022
rect 242164 177958 242216 177964
rect 240874 177576 240930 177585
rect 240874 177511 240930 177520
rect 242268 176225 242296 189790
rect 244936 176361 244964 302398
rect 246316 191350 246344 306410
rect 247684 295520 247736 295526
rect 247684 295462 247736 295468
rect 246396 254040 246448 254046
rect 246396 253982 246448 253988
rect 246304 191344 246356 191350
rect 246304 191286 246356 191292
rect 244922 176352 244978 176361
rect 244922 176287 244978 176296
rect 242254 176216 242310 176225
rect 239496 176180 239548 176186
rect 242254 176151 242310 176160
rect 239496 176122 239548 176128
rect 246408 176118 246436 253982
rect 247696 177614 247724 295462
rect 262220 294092 262272 294098
rect 262220 294034 262272 294040
rect 249064 291848 249116 291854
rect 249064 291790 249116 291796
rect 247776 280220 247828 280226
rect 247776 280162 247828 280168
rect 247788 194070 247816 280162
rect 247776 194064 247828 194070
rect 247776 194006 247828 194012
rect 249076 180794 249104 291790
rect 249156 291304 249208 291310
rect 249156 291246 249208 291252
rect 249168 189786 249196 291246
rect 251824 289876 251876 289882
rect 251824 289818 251876 289824
rect 249800 241528 249852 241534
rect 249800 241470 249852 241476
rect 249156 189780 249208 189786
rect 249156 189722 249208 189728
rect 249076 180766 249196 180794
rect 247684 177608 247736 177614
rect 247684 177550 247736 177556
rect 249064 176180 249116 176186
rect 249064 176122 249116 176128
rect 246396 176112 246448 176118
rect 246396 176054 246448 176060
rect 236644 175976 236696 175982
rect 236644 175918 236696 175924
rect 249076 172802 249104 176122
rect 249168 174321 249196 180766
rect 249340 178832 249392 178838
rect 249340 178774 249392 178780
rect 249248 176248 249300 176254
rect 249248 176190 249300 176196
rect 249260 175273 249288 176190
rect 249246 175264 249302 175273
rect 249246 175199 249302 175208
rect 249154 174312 249210 174321
rect 249154 174247 249210 174256
rect 249154 172816 249210 172825
rect 249076 172774 249154 172802
rect 249154 172751 249210 172760
rect 249352 172417 249380 178774
rect 249338 172408 249394 172417
rect 249338 172343 249394 172352
rect 249812 166705 249840 241470
rect 251836 198218 251864 289818
rect 255320 279472 255372 279478
rect 255320 279414 255372 279420
rect 252652 270564 252704 270570
rect 252652 270506 252704 270512
rect 252560 268388 252612 268394
rect 252560 268330 252612 268336
rect 251824 198212 251876 198218
rect 251824 198154 251876 198160
rect 251180 196716 251232 196722
rect 251180 196658 251232 196664
rect 249892 178016 249944 178022
rect 249892 177958 249944 177964
rect 249798 166696 249854 166705
rect 249798 166631 249854 166640
rect 249904 153513 249932 177958
rect 250626 159352 250682 159361
rect 250626 159287 250682 159296
rect 249890 153504 249946 153513
rect 249890 153439 249946 153448
rect 250444 138032 250496 138038
rect 250444 137974 250496 137980
rect 249154 96656 249210 96665
rect 249154 96591 249210 96600
rect 249064 95260 249116 95266
rect 249064 95202 249116 95208
rect 238024 93152 238076 93158
rect 238024 93094 238076 93100
rect 217324 3664 217376 3670
rect 217324 3606 217376 3612
rect 215944 3528 215996 3534
rect 215944 3470 215996 3476
rect 178684 3460 178736 3466
rect 178684 3402 178736 3408
rect 204904 3460 204956 3466
rect 204904 3402 204956 3408
rect 238036 2990 238064 93094
rect 249076 68338 249104 95202
rect 249064 68332 249116 68338
rect 249064 68274 249116 68280
rect 249168 34474 249196 96591
rect 249156 34468 249208 34474
rect 249156 34410 249208 34416
rect 248418 26888 248474 26897
rect 248418 26823 248474 26832
rect 244280 24268 244332 24274
rect 244280 24210 244332 24216
rect 241520 18760 241572 18766
rect 241520 18702 241572 18708
rect 241532 16574 241560 18702
rect 242992 17400 243044 17406
rect 242992 17342 243044 17348
rect 243004 16574 243032 17342
rect 244292 16574 244320 24210
rect 241532 16546 241744 16574
rect 243004 16546 244136 16574
rect 244292 16546 245240 16574
rect 239312 7744 239364 7750
rect 239312 7686 239364 7692
rect 235816 2984 235868 2990
rect 235816 2926 235868 2932
rect 238024 2984 238076 2990
rect 238024 2926 238076 2932
rect 235828 480 235856 2926
rect 239324 480 239352 7686
rect 240508 3596 240560 3602
rect 240508 3538 240560 3544
rect 240520 480 240548 3538
rect 241716 480 241744 16546
rect 242900 3664 242952 3670
rect 242900 3606 242952 3612
rect 242912 480 242940 3606
rect 244108 480 244136 16546
rect 245212 480 245240 16546
rect 247592 11892 247644 11898
rect 247592 11834 247644 11840
rect 246396 3460 246448 3466
rect 246396 3402 246448 3408
rect 246408 480 246436 3402
rect 247604 480 247632 11834
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 354 248460 26823
rect 250456 25702 250484 137974
rect 250536 136672 250588 136678
rect 250640 136649 250668 159287
rect 251192 157865 251220 196658
rect 251272 184340 251324 184346
rect 251272 184282 251324 184288
rect 251284 159633 251312 184282
rect 251364 178764 251416 178770
rect 251364 178706 251416 178712
rect 251376 171134 251404 178706
rect 252468 173868 252520 173874
rect 252468 173810 252520 173816
rect 252480 173777 252508 173810
rect 252466 173768 252522 173777
rect 252466 173703 252522 173712
rect 252468 172372 252520 172378
rect 252468 172314 252520 172320
rect 252480 171465 252508 172314
rect 252466 171456 252522 171465
rect 252466 171391 252522 171400
rect 251376 171106 251496 171134
rect 251364 165436 251416 165442
rect 251364 165378 251416 165384
rect 251376 164393 251404 165378
rect 251362 164384 251418 164393
rect 251362 164319 251418 164328
rect 251270 159624 251326 159633
rect 251270 159559 251326 159568
rect 251468 158817 251496 171106
rect 252376 171080 252428 171086
rect 252376 171022 252428 171028
rect 252284 170876 252336 170882
rect 252284 170818 252336 170824
rect 252296 170513 252324 170818
rect 252282 170504 252338 170513
rect 252282 170439 252338 170448
rect 252388 170105 252416 171022
rect 252466 170912 252522 170921
rect 252466 170847 252522 170856
rect 252480 170814 252508 170847
rect 252468 170808 252520 170814
rect 252468 170750 252520 170756
rect 252374 170096 252430 170105
rect 252374 170031 252430 170040
rect 252376 169720 252428 169726
rect 252376 169662 252428 169668
rect 252388 169153 252416 169662
rect 252466 169552 252522 169561
rect 252466 169487 252522 169496
rect 252374 169144 252430 169153
rect 252480 169114 252508 169487
rect 252374 169079 252430 169088
rect 252468 169108 252520 169114
rect 252468 169050 252520 169056
rect 252468 168700 252520 168706
rect 252468 168642 252520 168648
rect 252480 168609 252508 168642
rect 252466 168600 252522 168609
rect 252466 168535 252522 168544
rect 252376 168360 252428 168366
rect 252376 168302 252428 168308
rect 252388 167249 252416 168302
rect 252468 168292 252520 168298
rect 252468 168234 252520 168240
rect 252480 168201 252508 168234
rect 252466 168192 252522 168201
rect 252466 168127 252522 168136
rect 252466 167648 252522 167657
rect 252466 167583 252522 167592
rect 252480 167278 252508 167583
rect 252468 167272 252520 167278
rect 252374 167240 252430 167249
rect 252468 167214 252520 167220
rect 252374 167175 252430 167184
rect 252376 167000 252428 167006
rect 252376 166942 252428 166948
rect 252388 165753 252416 166942
rect 252468 166864 252520 166870
rect 252468 166806 252520 166812
rect 252480 166297 252508 166806
rect 252466 166288 252522 166297
rect 252466 166223 252522 166232
rect 252374 165744 252430 165753
rect 252374 165679 252430 165688
rect 252376 165572 252428 165578
rect 252376 165514 252428 165520
rect 252388 164801 252416 165514
rect 252468 165504 252520 165510
rect 252468 165446 252520 165452
rect 252480 165345 252508 165446
rect 252466 165336 252522 165345
rect 252466 165271 252522 165280
rect 252374 164792 252430 164801
rect 252374 164727 252430 164736
rect 252376 164212 252428 164218
rect 252376 164154 252428 164160
rect 252284 164144 252336 164150
rect 252284 164086 252336 164092
rect 252296 163033 252324 164086
rect 252388 163985 252416 164154
rect 252468 164076 252520 164082
rect 252468 164018 252520 164024
rect 252374 163976 252430 163985
rect 252374 163911 252430 163920
rect 252480 163441 252508 164018
rect 252466 163432 252522 163441
rect 252466 163367 252522 163376
rect 252282 163024 252338 163033
rect 252282 162959 252338 162968
rect 252468 162784 252520 162790
rect 252468 162726 252520 162732
rect 252480 161537 252508 162726
rect 252572 162489 252600 268330
rect 252664 171873 252692 270506
rect 253940 216028 253992 216034
rect 253940 215970 253992 215976
rect 252836 207732 252888 207738
rect 252836 207674 252888 207680
rect 252744 202224 252796 202230
rect 252744 202166 252796 202172
rect 252650 171864 252706 171873
rect 252650 171799 252706 171808
rect 252558 162480 252614 162489
rect 252558 162415 252614 162424
rect 252466 161528 252522 161537
rect 252466 161463 252522 161472
rect 252376 161424 252428 161430
rect 252376 161366 252428 161372
rect 252008 161016 252060 161022
rect 252008 160958 252060 160964
rect 252020 160177 252048 160958
rect 252388 160585 252416 161366
rect 252466 161120 252522 161129
rect 252466 161055 252522 161064
rect 252480 160818 252508 161055
rect 252468 160812 252520 160818
rect 252468 160754 252520 160760
rect 252374 160576 252430 160585
rect 252374 160511 252430 160520
rect 252006 160168 252062 160177
rect 252006 160103 252062 160112
rect 252468 160064 252520 160070
rect 252468 160006 252520 160012
rect 252480 159225 252508 160006
rect 252466 159216 252522 159225
rect 252466 159151 252522 159160
rect 251454 158808 251510 158817
rect 251454 158743 251510 158752
rect 252468 158704 252520 158710
rect 252006 158672 252062 158681
rect 252468 158646 252520 158652
rect 252006 158607 252062 158616
rect 251178 157856 251234 157865
rect 251178 157791 251234 157800
rect 251548 155848 251600 155854
rect 251548 155790 251600 155796
rect 251560 155417 251588 155790
rect 251546 155408 251602 155417
rect 251546 155343 251602 155352
rect 251824 153876 251876 153882
rect 251824 153818 251876 153824
rect 251364 151496 251416 151502
rect 251364 151438 251416 151444
rect 251376 150793 251404 151438
rect 251362 150784 251418 150793
rect 251362 150719 251418 150728
rect 251640 143404 251692 143410
rect 251640 143346 251692 143352
rect 251652 142769 251680 143346
rect 251638 142760 251694 142769
rect 251638 142695 251694 142704
rect 250536 136614 250588 136620
rect 250626 136640 250682 136649
rect 250548 49162 250576 136614
rect 250626 136575 250682 136584
rect 251732 126880 251784 126886
rect 251732 126822 251784 126828
rect 251744 125769 251772 126822
rect 251730 125760 251786 125769
rect 251730 125695 251786 125704
rect 251836 115433 251864 153818
rect 251916 140820 251968 140826
rect 251916 140762 251968 140768
rect 251822 115424 251878 115433
rect 251822 115359 251878 115368
rect 251928 114481 251956 140762
rect 252020 140457 252048 158607
rect 252480 158273 252508 158646
rect 252466 158264 252522 158273
rect 252466 158199 252522 158208
rect 252376 157344 252428 157350
rect 252376 157286 252428 157292
rect 252388 156369 252416 157286
rect 252468 157276 252520 157282
rect 252468 157218 252520 157224
rect 252480 156913 252508 157218
rect 252466 156904 252522 156913
rect 252466 156839 252522 156848
rect 252374 156360 252430 156369
rect 252374 156295 252430 156304
rect 252466 155952 252522 155961
rect 252466 155887 252468 155896
rect 252520 155887 252522 155896
rect 252468 155858 252520 155864
rect 252468 155780 252520 155786
rect 252468 155722 252520 155728
rect 252480 155009 252508 155722
rect 252466 155000 252522 155009
rect 252466 154935 252522 154944
rect 252468 154488 252520 154494
rect 252468 154430 252520 154436
rect 252480 154057 252508 154430
rect 252466 154048 252522 154057
rect 252466 153983 252522 153992
rect 252376 153196 252428 153202
rect 252376 153138 252428 153144
rect 252388 152697 252416 153138
rect 252468 153128 252520 153134
rect 252466 153096 252468 153105
rect 252520 153096 252522 153105
rect 252466 153031 252522 153040
rect 252374 152688 252430 152697
rect 252374 152623 252430 152632
rect 252468 151768 252520 151774
rect 252374 151736 252430 151745
rect 252468 151710 252520 151716
rect 252374 151671 252376 151680
rect 252428 151671 252430 151680
rect 252376 151642 252428 151648
rect 252480 151201 252508 151710
rect 252466 151192 252522 151201
rect 252466 151127 252522 151136
rect 252468 150408 252520 150414
rect 252468 150350 252520 150356
rect 252100 150340 252152 150346
rect 252100 150282 252152 150288
rect 252112 149841 252140 150282
rect 252284 150272 252336 150278
rect 252480 150249 252508 150350
rect 252284 150214 252336 150220
rect 252466 150240 252522 150249
rect 252098 149832 252154 149841
rect 252098 149767 252154 149776
rect 252296 149297 252324 150214
rect 252466 150175 252522 150184
rect 252282 149288 252338 149297
rect 252282 149223 252338 149232
rect 252376 149048 252428 149054
rect 252376 148990 252428 148996
rect 252284 148912 252336 148918
rect 252284 148854 252336 148860
rect 252296 147937 252324 148854
rect 252388 148345 252416 148990
rect 252468 148980 252520 148986
rect 252468 148922 252520 148928
rect 252480 148889 252508 148922
rect 252466 148880 252522 148889
rect 252466 148815 252522 148824
rect 252374 148336 252430 148345
rect 252374 148271 252430 148280
rect 252282 147928 252338 147937
rect 252282 147863 252338 147872
rect 252468 147552 252520 147558
rect 252468 147494 252520 147500
rect 252192 146940 252244 146946
rect 252192 146882 252244 146888
rect 252204 144673 252232 146882
rect 252480 146577 252508 147494
rect 252756 146985 252784 202166
rect 252848 154465 252876 207674
rect 252834 154456 252890 154465
rect 252834 154391 252890 154400
rect 253952 151502 253980 215970
rect 254124 213376 254176 213382
rect 254124 213318 254176 213324
rect 254032 209228 254084 209234
rect 254032 209170 254084 209176
rect 254044 155922 254072 209170
rect 254136 165442 254164 213318
rect 254216 192568 254268 192574
rect 254216 192510 254268 192516
rect 254124 165436 254176 165442
rect 254124 165378 254176 165384
rect 254032 155916 254084 155922
rect 254032 155858 254084 155864
rect 254228 155854 254256 192510
rect 255332 161022 255360 279414
rect 256976 218816 257028 218822
rect 256976 218758 257028 218764
rect 255412 206304 255464 206310
rect 255412 206246 255464 206252
rect 255320 161016 255372 161022
rect 255320 160958 255372 160964
rect 254584 158772 254636 158778
rect 254584 158714 254636 158720
rect 254216 155848 254268 155854
rect 254216 155790 254268 155796
rect 253940 151496 253992 151502
rect 253940 151438 253992 151444
rect 252742 146976 252798 146985
rect 252742 146911 252798 146920
rect 252466 146568 252522 146577
rect 252466 146503 252522 146512
rect 252468 146260 252520 146266
rect 252468 146202 252520 146208
rect 252376 146192 252428 146198
rect 252376 146134 252428 146140
rect 252284 146124 252336 146130
rect 252284 146066 252336 146072
rect 252296 145081 252324 146066
rect 252388 145625 252416 146134
rect 252480 146033 252508 146202
rect 252466 146024 252522 146033
rect 252466 145959 252522 145968
rect 252374 145616 252430 145625
rect 252374 145551 252430 145560
rect 253480 145580 253532 145586
rect 253480 145522 253532 145528
rect 252282 145072 252338 145081
rect 252282 145007 252338 145016
rect 252376 144900 252428 144906
rect 252376 144842 252428 144848
rect 252190 144664 252246 144673
rect 252190 144599 252246 144608
rect 252388 143721 252416 144842
rect 252468 144832 252520 144838
rect 252468 144774 252520 144780
rect 252480 144129 252508 144774
rect 253388 144220 253440 144226
rect 253388 144162 253440 144168
rect 252466 144120 252522 144129
rect 252466 144055 252522 144064
rect 252374 143712 252430 143721
rect 252374 143647 252430 143656
rect 252376 143540 252428 143546
rect 252376 143482 252428 143488
rect 252388 142225 252416 143482
rect 252468 143472 252520 143478
rect 252468 143414 252520 143420
rect 252480 143177 252508 143414
rect 252466 143168 252522 143177
rect 252466 143103 252522 143112
rect 252374 142216 252430 142225
rect 252374 142151 252430 142160
rect 253296 142180 253348 142186
rect 253296 142122 253348 142128
rect 252376 142112 252428 142118
rect 252376 142054 252428 142060
rect 252388 140865 252416 142054
rect 253202 141672 253258 141681
rect 253202 141607 253258 141616
rect 252466 141400 252522 141409
rect 252466 141335 252522 141344
rect 252480 141166 252508 141335
rect 252468 141160 252520 141166
rect 252468 141102 252520 141108
rect 252374 140856 252430 140865
rect 252374 140791 252430 140800
rect 252468 140752 252520 140758
rect 252468 140694 252520 140700
rect 252376 140684 252428 140690
rect 252376 140626 252428 140632
rect 252006 140448 252062 140457
rect 252006 140383 252062 140392
rect 252100 140072 252152 140078
rect 252100 140014 252152 140020
rect 252008 136400 252060 136406
rect 252008 136342 252060 136348
rect 252020 118833 252048 136342
rect 252112 129169 252140 140014
rect 252388 139505 252416 140626
rect 252480 139913 252508 140694
rect 252466 139904 252522 139913
rect 252466 139839 252522 139848
rect 252374 139496 252430 139505
rect 252374 139431 252430 139440
rect 252376 139392 252428 139398
rect 252376 139334 252428 139340
rect 252388 138553 252416 139334
rect 252468 139324 252520 139330
rect 252468 139266 252520 139272
rect 252480 138961 252508 139266
rect 252466 138952 252522 138961
rect 252466 138887 252522 138896
rect 252374 138544 252430 138553
rect 252374 138479 252430 138488
rect 252468 137964 252520 137970
rect 252468 137906 252520 137912
rect 252376 137896 252428 137902
rect 252376 137838 252428 137844
rect 252388 137057 252416 137838
rect 252480 137601 252508 137906
rect 252466 137592 252522 137601
rect 252466 137527 252522 137536
rect 252374 137048 252430 137057
rect 252374 136983 252430 136992
rect 252284 136604 252336 136610
rect 252284 136546 252336 136552
rect 252296 135289 252324 136546
rect 252468 136536 252520 136542
rect 252468 136478 252520 136484
rect 252376 136468 252428 136474
rect 252376 136410 252428 136416
rect 252388 135697 252416 136410
rect 252480 136241 252508 136478
rect 252466 136232 252522 136241
rect 252466 136167 252522 136176
rect 252374 135688 252430 135697
rect 252374 135623 252430 135632
rect 252282 135280 252338 135289
rect 252282 135215 252338 135224
rect 252376 135244 252428 135250
rect 252376 135186 252428 135192
rect 252388 134337 252416 135186
rect 252468 135176 252520 135182
rect 252468 135118 252520 135124
rect 252480 134745 252508 135118
rect 252466 134736 252522 134745
rect 252466 134671 252522 134680
rect 252374 134328 252430 134337
rect 252374 134263 252430 134272
rect 252376 133884 252428 133890
rect 252376 133826 252428 133832
rect 252284 133816 252336 133822
rect 252284 133758 252336 133764
rect 252296 132841 252324 133758
rect 252388 133385 252416 133826
rect 252466 133784 252522 133793
rect 252466 133719 252468 133728
rect 252520 133719 252522 133728
rect 252468 133690 252520 133696
rect 252374 133376 252430 133385
rect 252374 133311 252430 133320
rect 252282 132832 252338 132841
rect 252282 132767 252338 132776
rect 252284 132456 252336 132462
rect 252284 132398 252336 132404
rect 252466 132424 252522 132433
rect 252296 131481 252324 132398
rect 252376 132388 252428 132394
rect 252466 132359 252522 132368
rect 252376 132330 252428 132336
rect 252388 131889 252416 132330
rect 252480 132326 252508 132359
rect 252468 132320 252520 132326
rect 252468 132262 252520 132268
rect 252374 131880 252430 131889
rect 252374 131815 252430 131824
rect 252282 131472 252338 131481
rect 252282 131407 252338 131416
rect 252468 131096 252520 131102
rect 252468 131038 252520 131044
rect 252376 131028 252428 131034
rect 252376 130970 252428 130976
rect 252284 130960 252336 130966
rect 252284 130902 252336 130908
rect 252296 130121 252324 130902
rect 252388 130529 252416 130970
rect 252480 130937 252508 131038
rect 252466 130928 252522 130937
rect 252466 130863 252522 130872
rect 252374 130520 252430 130529
rect 252374 130455 252430 130464
rect 252282 130112 252338 130121
rect 252282 130047 252338 130056
rect 252376 129736 252428 129742
rect 252376 129678 252428 129684
rect 252098 129160 252154 129169
rect 252098 129095 252154 129104
rect 252388 128625 252416 129678
rect 252468 129668 252520 129674
rect 252468 129610 252520 129616
rect 252480 129577 252508 129610
rect 252466 129568 252522 129577
rect 252466 129503 252522 129512
rect 252374 128616 252430 128625
rect 252374 128551 252430 128560
rect 252192 128376 252244 128382
rect 252192 128318 252244 128324
rect 252204 126313 252232 128318
rect 252468 128308 252520 128314
rect 252468 128250 252520 128256
rect 252284 128240 252336 128246
rect 252480 128217 252508 128250
rect 252284 128182 252336 128188
rect 252466 128208 252522 128217
rect 252296 127673 252324 128182
rect 252376 128172 252428 128178
rect 252466 128143 252522 128152
rect 252376 128114 252428 128120
rect 252282 127664 252338 127673
rect 252282 127599 252338 127608
rect 252388 127265 252416 128114
rect 252374 127256 252430 127265
rect 252374 127191 252430 127200
rect 252468 126948 252520 126954
rect 252468 126890 252520 126896
rect 252480 126721 252508 126890
rect 252466 126712 252522 126721
rect 252466 126647 252522 126656
rect 252190 126304 252246 126313
rect 252190 126239 252246 126248
rect 252284 126268 252336 126274
rect 252284 126210 252336 126216
rect 252296 125361 252324 126210
rect 252468 125588 252520 125594
rect 252468 125530 252520 125536
rect 252376 125520 252428 125526
rect 252376 125462 252428 125468
rect 252282 125352 252338 125361
rect 252282 125287 252338 125296
rect 252388 124409 252416 125462
rect 252480 124817 252508 125530
rect 252466 124808 252522 124817
rect 252466 124743 252522 124752
rect 252374 124400 252430 124409
rect 252374 124335 252430 124344
rect 252468 124160 252520 124166
rect 252468 124102 252520 124108
rect 252376 124092 252428 124098
rect 252376 124034 252428 124040
rect 252284 124024 252336 124030
rect 252284 123966 252336 123972
rect 252296 123049 252324 123966
rect 252388 123457 252416 124034
rect 252480 124001 252508 124102
rect 252466 123992 252522 124001
rect 252466 123927 252522 123936
rect 252374 123448 252430 123457
rect 252374 123383 252430 123392
rect 252282 123040 252338 123049
rect 252282 122975 252338 122984
rect 252468 122800 252520 122806
rect 252468 122742 252520 122748
rect 252284 122732 252336 122738
rect 252284 122674 252336 122680
rect 252296 122097 252324 122674
rect 252480 122505 252508 122742
rect 252466 122496 252522 122505
rect 252376 122460 252428 122466
rect 252466 122431 252522 122440
rect 252376 122402 252428 122408
rect 252282 122088 252338 122097
rect 252282 122023 252338 122032
rect 252388 121553 252416 122402
rect 252374 121544 252430 121553
rect 252374 121479 252430 121488
rect 252376 121440 252428 121446
rect 252376 121382 252428 121388
rect 252388 120601 252416 121382
rect 252468 121372 252520 121378
rect 252468 121314 252520 121320
rect 252480 121145 252508 121314
rect 252466 121136 252522 121145
rect 252466 121071 252522 121080
rect 252468 120964 252520 120970
rect 252468 120906 252520 120912
rect 252374 120592 252430 120601
rect 252374 120527 252430 120536
rect 252480 120193 252508 120906
rect 252466 120184 252522 120193
rect 252466 120119 252522 120128
rect 252468 120080 252520 120086
rect 252468 120022 252520 120028
rect 252284 120012 252336 120018
rect 252284 119954 252336 119960
rect 252296 119241 252324 119954
rect 252480 119649 252508 120022
rect 252466 119640 252522 119649
rect 252466 119575 252522 119584
rect 252376 119400 252428 119406
rect 252376 119342 252428 119348
rect 252282 119232 252338 119241
rect 252282 119167 252338 119176
rect 252006 118824 252062 118833
rect 252006 118759 252062 118768
rect 252388 117337 252416 119342
rect 252468 118652 252520 118658
rect 252468 118594 252520 118600
rect 252480 118289 252508 118594
rect 252466 118280 252522 118289
rect 252466 118215 252522 118224
rect 252466 117872 252522 117881
rect 252466 117807 252522 117816
rect 252480 117706 252508 117807
rect 252468 117700 252520 117706
rect 252468 117642 252520 117648
rect 252374 117328 252430 117337
rect 252374 117263 252430 117272
rect 252468 117292 252520 117298
rect 252468 117234 252520 117240
rect 252376 117224 252428 117230
rect 252376 117166 252428 117172
rect 252388 116385 252416 117166
rect 252480 116929 252508 117234
rect 252466 116920 252522 116929
rect 252466 116855 252522 116864
rect 252468 116544 252520 116550
rect 252468 116486 252520 116492
rect 252374 116376 252430 116385
rect 252374 116311 252430 116320
rect 252480 115977 252508 116486
rect 252466 115968 252522 115977
rect 252376 115932 252428 115938
rect 252466 115903 252522 115912
rect 252376 115874 252428 115880
rect 252388 115025 252416 115874
rect 252468 115252 252520 115258
rect 252468 115194 252520 115200
rect 252374 115016 252430 115025
rect 252374 114951 252430 114960
rect 252480 114594 252508 115194
rect 252388 114566 252508 114594
rect 251914 114472 251970 114481
rect 251914 114407 251970 114416
rect 252284 114436 252336 114442
rect 252284 114378 252336 114384
rect 251732 114368 251784 114374
rect 251732 114310 251784 114316
rect 251744 113529 251772 114310
rect 251730 113520 251786 113529
rect 251730 113455 251786 113464
rect 252100 112464 252152 112470
rect 252100 112406 252152 112412
rect 251732 108860 251784 108866
rect 251732 108802 251784 108808
rect 251744 108361 251772 108802
rect 251730 108352 251786 108361
rect 251730 108287 251786 108296
rect 251180 106208 251232 106214
rect 251180 106150 251232 106156
rect 251192 106049 251220 106150
rect 251178 106040 251234 106049
rect 251178 105975 251234 105984
rect 252112 103737 252140 112406
rect 252296 111217 252324 114378
rect 252388 112713 252416 114566
rect 252468 114504 252520 114510
rect 252468 114446 252520 114452
rect 252480 114073 252508 114446
rect 252466 114064 252522 114073
rect 252466 113999 252522 114008
rect 252468 113144 252520 113150
rect 252466 113112 252468 113121
rect 252520 113112 252522 113121
rect 252466 113047 252522 113056
rect 252374 112704 252430 112713
rect 252374 112639 252430 112648
rect 252468 112328 252520 112334
rect 252468 112270 252520 112276
rect 252480 112169 252508 112270
rect 252466 112160 252522 112169
rect 252466 112095 252522 112104
rect 252468 111784 252520 111790
rect 252466 111752 252468 111761
rect 252520 111752 252522 111761
rect 252376 111716 252428 111722
rect 252466 111687 252522 111696
rect 252376 111658 252428 111664
rect 252282 111208 252338 111217
rect 252282 111143 252338 111152
rect 252388 110809 252416 111658
rect 252374 110800 252430 110809
rect 252374 110735 252430 110744
rect 252192 110560 252244 110566
rect 252192 110502 252244 110508
rect 252204 105097 252232 110502
rect 252376 110424 252428 110430
rect 252376 110366 252428 110372
rect 252284 110288 252336 110294
rect 252284 110230 252336 110236
rect 252296 109313 252324 110230
rect 252388 109857 252416 110366
rect 252468 110356 252520 110362
rect 252468 110298 252520 110304
rect 252480 110265 252508 110298
rect 252466 110256 252522 110265
rect 252466 110191 252522 110200
rect 252374 109848 252430 109857
rect 252374 109783 252430 109792
rect 252282 109304 252338 109313
rect 252282 109239 252338 109248
rect 252376 108996 252428 109002
rect 252376 108938 252428 108944
rect 252388 107953 252416 108938
rect 252468 108928 252520 108934
rect 252466 108896 252468 108905
rect 252520 108896 252522 108905
rect 252466 108831 252522 108840
rect 252374 107944 252430 107953
rect 252374 107879 252430 107888
rect 252376 107636 252428 107642
rect 252376 107578 252428 107584
rect 252284 107500 252336 107506
rect 252284 107442 252336 107448
rect 252296 107001 252324 107442
rect 252282 106992 252338 107001
rect 252282 106927 252338 106936
rect 252388 106593 252416 107578
rect 252468 107568 252520 107574
rect 252466 107536 252468 107545
rect 252520 107536 252522 107545
rect 252466 107471 252522 107480
rect 252374 106584 252430 106593
rect 252374 106519 252430 106528
rect 252468 106276 252520 106282
rect 252468 106218 252520 106224
rect 252480 105641 252508 106218
rect 252466 105632 252522 105641
rect 252466 105567 252522 105576
rect 252376 105528 252428 105534
rect 252376 105470 252428 105476
rect 252190 105088 252246 105097
rect 252190 105023 252246 105032
rect 252098 103728 252154 103737
rect 252098 103663 252154 103672
rect 252284 103216 252336 103222
rect 252284 103158 252336 103164
rect 252192 103148 252244 103154
rect 252192 103090 252244 103096
rect 252204 102785 252232 103090
rect 252190 102776 252246 102785
rect 252190 102711 252246 102720
rect 252192 101448 252244 101454
rect 252296 101425 252324 103158
rect 252388 102241 252416 105470
rect 252468 104848 252520 104854
rect 252468 104790 252520 104796
rect 252480 104145 252508 104790
rect 252466 104136 252522 104145
rect 252466 104071 252522 104080
rect 252468 104032 252520 104038
rect 252468 103974 252520 103980
rect 252480 103193 252508 103974
rect 252466 103184 252522 103193
rect 252466 103119 252522 103128
rect 252374 102232 252430 102241
rect 252374 102167 252430 102176
rect 252468 102128 252520 102134
rect 252468 102070 252520 102076
rect 252192 101390 252244 101396
rect 252282 101416 252338 101425
rect 252204 97617 252232 101390
rect 252282 101351 252338 101360
rect 252480 100881 252508 102070
rect 252466 100872 252522 100881
rect 252466 100807 252522 100816
rect 252284 100700 252336 100706
rect 252284 100642 252336 100648
rect 252296 99521 252324 100642
rect 252468 100632 252520 100638
rect 252468 100574 252520 100580
rect 252376 100564 252428 100570
rect 252376 100506 252428 100512
rect 252388 99929 252416 100506
rect 252480 100473 252508 100574
rect 252466 100464 252522 100473
rect 252466 100399 252522 100408
rect 252374 99920 252430 99929
rect 252374 99855 252430 99864
rect 252282 99512 252338 99521
rect 252282 99447 252338 99456
rect 252468 99272 252520 99278
rect 252468 99214 252520 99220
rect 252376 99204 252428 99210
rect 252376 99146 252428 99152
rect 252388 98025 252416 99146
rect 252480 98569 252508 99214
rect 253216 98977 253244 141607
rect 253308 103222 253336 142122
rect 253400 106214 253428 144162
rect 253492 120018 253520 145522
rect 254596 136406 254624 158714
rect 254860 154624 254912 154630
rect 254860 154566 254912 154572
rect 254768 153264 254820 153270
rect 254768 153206 254820 153212
rect 254676 149116 254728 149122
rect 254676 149058 254728 149064
rect 254584 136400 254636 136406
rect 254584 136342 254636 136348
rect 254584 125656 254636 125662
rect 254584 125598 254636 125604
rect 253480 120012 253532 120018
rect 253480 119954 253532 119960
rect 253388 106208 253440 106214
rect 253388 106150 253440 106156
rect 253296 103216 253348 103222
rect 253296 103158 253348 103164
rect 253388 102196 253440 102202
rect 253388 102138 253440 102144
rect 253202 98968 253258 98977
rect 253202 98903 253258 98912
rect 252466 98560 252522 98569
rect 252466 98495 252522 98504
rect 252374 98016 252430 98025
rect 252374 97951 252430 97960
rect 252190 97608 252246 97617
rect 252190 97543 252246 97552
rect 252468 97300 252520 97306
rect 252468 97242 252520 97248
rect 252480 97073 252508 97242
rect 251270 97064 251326 97073
rect 251270 96999 251326 97008
rect 252466 97064 252522 97073
rect 252466 96999 252522 97008
rect 251178 96248 251234 96257
rect 251178 96183 251234 96192
rect 251192 93922 251220 96183
rect 251100 93894 251220 93922
rect 251100 93854 251128 93894
rect 251100 93826 251220 93854
rect 251192 93158 251220 93826
rect 251180 93152 251232 93158
rect 251180 93094 251232 93100
rect 251284 84194 251312 96999
rect 253204 96688 253256 96694
rect 253204 96630 253256 96636
rect 251192 84166 251312 84194
rect 250536 49156 250588 49162
rect 250536 49098 250588 49104
rect 251192 35902 251220 84166
rect 251180 35896 251232 35902
rect 251180 35838 251232 35844
rect 251180 29776 251232 29782
rect 251180 29718 251232 29724
rect 250444 25696 250496 25702
rect 250444 25638 250496 25644
rect 249984 7676 250036 7682
rect 249984 7618 250036 7624
rect 249996 480 250024 7618
rect 251192 3602 251220 29718
rect 253216 29714 253244 96630
rect 253400 71058 253428 102138
rect 254596 73982 254624 125598
rect 254688 108866 254716 149058
rect 254780 114374 254808 153206
rect 254872 140826 254900 154566
rect 255424 151706 255452 206246
rect 255504 200932 255556 200938
rect 255504 200874 255556 200880
rect 255412 151700 255464 151706
rect 255412 151642 255464 151648
rect 255516 150346 255544 200874
rect 256792 191208 256844 191214
rect 256792 191150 256844 191156
rect 255596 176112 255648 176118
rect 255596 176054 255648 176060
rect 255504 150340 255556 150346
rect 255504 150282 255556 150288
rect 255608 150278 255636 176054
rect 256148 151836 256200 151842
rect 256148 151778 256200 151784
rect 256056 150476 256108 150482
rect 256056 150418 256108 150424
rect 255596 150272 255648 150278
rect 255596 150214 255648 150220
rect 255320 149388 255372 149394
rect 255320 149330 255372 149336
rect 255332 143410 255360 149330
rect 255320 143404 255372 143410
rect 255320 143346 255372 143352
rect 254860 140820 254912 140826
rect 254860 140762 254912 140768
rect 254860 137284 254912 137290
rect 254860 137226 254912 137232
rect 254872 126886 254900 137226
rect 254860 126880 254912 126886
rect 254860 126822 254912 126828
rect 255964 124228 256016 124234
rect 255964 124170 256016 124176
rect 254768 114368 254820 114374
rect 254768 114310 254820 114316
rect 254676 108860 254728 108866
rect 254676 108802 254728 108808
rect 255318 80744 255374 80753
rect 255318 80679 255374 80688
rect 254584 73976 254636 73982
rect 254584 73918 254636 73924
rect 253388 71052 253440 71058
rect 253388 70994 253440 71000
rect 253204 29708 253256 29714
rect 253204 29650 253256 29656
rect 255332 16574 255360 80679
rect 255976 72622 256004 124170
rect 256068 110294 256096 150418
rect 256160 114442 256188 151778
rect 256804 148918 256832 191150
rect 256884 175976 256936 175982
rect 256884 175918 256936 175924
rect 256896 170882 256924 175918
rect 256884 170876 256936 170882
rect 256884 170818 256936 170824
rect 256792 148912 256844 148918
rect 256792 148854 256844 148860
rect 256240 146328 256292 146334
rect 256240 146270 256292 146276
rect 256148 114436 256200 114442
rect 256148 114378 256200 114384
rect 256252 110566 256280 146270
rect 256988 140690 257016 218758
rect 259460 204944 259512 204950
rect 259460 204886 259512 204892
rect 258264 183184 258316 183190
rect 258264 183126 258316 183132
rect 258080 181756 258132 181762
rect 258080 181698 258132 181704
rect 257528 162920 257580 162926
rect 257528 162862 257580 162868
rect 257344 147824 257396 147830
rect 257344 147766 257396 147772
rect 256976 140684 257028 140690
rect 256976 140626 257028 140632
rect 256240 110560 256292 110566
rect 256240 110502 256292 110508
rect 256056 110288 256108 110294
rect 256056 110230 256108 110236
rect 257356 107506 257384 147766
rect 257436 143608 257488 143614
rect 257436 143550 257488 143556
rect 257344 107500 257396 107506
rect 257344 107442 257396 107448
rect 257448 103154 257476 143550
rect 257540 124030 257568 162862
rect 258092 149394 258120 181698
rect 258172 177608 258224 177614
rect 258172 177550 258224 177556
rect 258184 160818 258212 177550
rect 258276 170814 258304 183126
rect 258356 180464 258408 180470
rect 258356 180406 258408 180412
rect 258264 170808 258316 170814
rect 258264 170750 258316 170756
rect 258368 169114 258396 180406
rect 259092 169788 259144 169794
rect 259092 169730 259144 169736
rect 258356 169108 258408 169114
rect 258356 169050 258408 169056
rect 259104 167278 259132 169730
rect 259092 167272 259144 167278
rect 259092 167214 259144 167220
rect 259472 166870 259500 204886
rect 260840 200864 260892 200870
rect 260840 200806 260892 200812
rect 259736 193996 259788 194002
rect 259736 193938 259788 193944
rect 259552 178900 259604 178906
rect 259552 178842 259604 178848
rect 259460 166864 259512 166870
rect 259460 166806 259512 166812
rect 258908 161492 258960 161498
rect 258908 161434 258960 161440
rect 258172 160812 258224 160818
rect 258172 160754 258224 160760
rect 258724 160132 258776 160138
rect 258724 160074 258776 160080
rect 258080 149388 258132 149394
rect 258080 149330 258132 149336
rect 257528 124024 257580 124030
rect 257528 123966 257580 123972
rect 258736 120970 258764 160074
rect 258816 157412 258868 157418
rect 258816 157354 258868 157360
rect 258724 120964 258776 120970
rect 258724 120906 258776 120912
rect 258828 117706 258856 157354
rect 258920 122466 258948 161434
rect 259000 148368 259052 148374
rect 259000 148310 259052 148316
rect 258908 122460 258960 122466
rect 258908 122402 258960 122408
rect 258816 117700 258868 117706
rect 258816 117642 258868 117648
rect 259012 112334 259040 148310
rect 259564 141166 259592 178842
rect 259644 177472 259696 177478
rect 259644 177414 259696 177420
rect 259656 146130 259684 177414
rect 259748 168706 259776 193938
rect 260852 169726 260880 200806
rect 261024 196784 261076 196790
rect 261024 196726 261076 196732
rect 260932 177540 260984 177546
rect 260932 177482 260984 177488
rect 260840 169720 260892 169726
rect 260840 169662 260892 169668
rect 259736 168700 259788 168706
rect 259736 168642 259788 168648
rect 260196 165640 260248 165646
rect 260196 165582 260248 165588
rect 260104 155984 260156 155990
rect 260104 155926 260156 155932
rect 259644 146124 259696 146130
rect 259644 146066 259696 146072
rect 259552 141160 259604 141166
rect 259552 141102 259604 141108
rect 260116 116550 260144 155926
rect 260208 128382 260236 165582
rect 260944 146946 260972 177482
rect 261036 167006 261064 196726
rect 261116 188692 261168 188698
rect 261116 188634 261168 188640
rect 261024 167000 261076 167006
rect 261024 166942 261076 166948
rect 261128 165510 261156 188634
rect 262232 169794 262260 294034
rect 263600 252680 263652 252686
rect 263600 252622 263652 252628
rect 262312 191140 262364 191146
rect 262312 191082 262364 191088
rect 262220 169788 262272 169794
rect 262220 169730 262272 169736
rect 261116 165504 261168 165510
rect 261116 165446 261168 165452
rect 260932 146940 260984 146946
rect 260932 146882 260984 146888
rect 261484 146396 261536 146402
rect 261484 146338 261536 146344
rect 260196 128376 260248 128382
rect 260196 128318 260248 128324
rect 260104 116544 260156 116550
rect 260104 116486 260156 116492
rect 260104 113212 260156 113218
rect 260104 113154 260156 113160
rect 259000 112328 259052 112334
rect 259000 112270 259052 112276
rect 258724 105052 258776 105058
rect 258724 104994 258776 105000
rect 257436 103148 257488 103154
rect 257436 103090 257488 103096
rect 257344 102264 257396 102270
rect 257344 102206 257396 102212
rect 255964 72616 256016 72622
rect 255964 72558 256016 72564
rect 255332 16546 255912 16574
rect 251270 13152 251326 13161
rect 251270 13087 251326 13096
rect 251180 3596 251232 3602
rect 251180 3538 251232 3544
rect 251284 3482 251312 13087
rect 254676 9104 254728 9110
rect 254676 9046 254728 9052
rect 252376 3596 252428 3602
rect 252376 3538 252428 3544
rect 251192 3454 251312 3482
rect 251192 480 251220 3454
rect 252388 480 252416 3538
rect 253480 3528 253532 3534
rect 253480 3470 253532 3476
rect 253492 480 253520 3470
rect 254688 480 254716 9046
rect 255884 480 255912 16546
rect 257356 14550 257384 102206
rect 257344 14544 257396 14550
rect 257344 14486 257396 14492
rect 256700 10464 256752 10470
rect 256700 10406 256752 10412
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 256712 354 256740 10406
rect 258736 4826 258764 104994
rect 260116 50386 260144 113154
rect 261496 106282 261524 146338
rect 262324 139330 262352 191082
rect 262404 188556 262456 188562
rect 262404 188498 262456 188504
rect 262416 168298 262444 188498
rect 262496 177404 262548 177410
rect 262496 177346 262548 177352
rect 262404 168292 262456 168298
rect 262404 168234 262456 168240
rect 262508 144838 262536 177346
rect 262864 168428 262916 168434
rect 262864 168370 262916 168376
rect 262496 144832 262548 144838
rect 262496 144774 262548 144780
rect 262312 139324 262364 139330
rect 262312 139266 262364 139272
rect 262876 130966 262904 168370
rect 263612 168366 263640 252622
rect 266360 247104 266412 247110
rect 266360 247046 266412 247052
rect 263784 203584 263836 203590
rect 263784 203526 263836 203532
rect 263692 180328 263744 180334
rect 263692 180270 263744 180276
rect 263600 168360 263652 168366
rect 263600 168302 263652 168308
rect 262956 158840 263008 158846
rect 262956 158782 263008 158788
rect 262864 130960 262916 130966
rect 262864 130902 262916 130908
rect 262968 120086 262996 158782
rect 263704 143478 263732 180270
rect 263796 173874 263824 203526
rect 265072 199572 265124 199578
rect 265072 199514 265124 199520
rect 263876 183116 263928 183122
rect 263876 183058 263928 183064
rect 263784 173868 263836 173874
rect 263784 173810 263836 173816
rect 263888 164082 263916 183058
rect 264980 181688 265032 181694
rect 264980 181630 265032 181636
rect 264428 171148 264480 171154
rect 264428 171090 264480 171096
rect 263876 164076 263928 164082
rect 263876 164018 263928 164024
rect 264244 161560 264296 161566
rect 264244 161502 264296 161508
rect 263692 143472 263744 143478
rect 263692 143414 263744 143420
rect 264256 122738 264284 161502
rect 264336 157480 264388 157486
rect 264336 157422 264388 157428
rect 264244 122732 264296 122738
rect 264244 122674 264296 122680
rect 262956 120080 263008 120086
rect 262956 120022 263008 120028
rect 262864 118720 262916 118726
rect 262864 118662 262916 118668
rect 261484 106276 261536 106282
rect 261484 106218 261536 106224
rect 261484 98048 261536 98054
rect 261484 97990 261536 97996
rect 260840 78056 260892 78062
rect 260840 77998 260892 78004
rect 260104 50380 260156 50386
rect 260104 50322 260156 50328
rect 260852 16574 260880 77998
rect 261496 22778 261524 97990
rect 262876 46306 262904 118662
rect 264348 118658 264376 157422
rect 264440 132326 264468 171090
rect 264992 143546 265020 181630
rect 265084 171086 265112 199514
rect 265256 180396 265308 180402
rect 265256 180338 265308 180344
rect 265164 178968 265216 178974
rect 265164 178910 265216 178916
rect 265072 171080 265124 171086
rect 265072 171022 265124 171028
rect 265176 157282 265204 178910
rect 265268 164150 265296 180338
rect 266372 172378 266400 247046
rect 267740 231124 267792 231130
rect 267740 231066 267792 231072
rect 266452 185972 266504 185978
rect 266452 185914 266504 185920
rect 266360 172372 266412 172378
rect 266360 172314 266412 172320
rect 265256 164144 265308 164150
rect 265256 164086 265308 164092
rect 265624 160200 265676 160206
rect 265624 160142 265676 160148
rect 265164 157276 265216 157282
rect 265164 157218 265216 157224
rect 264980 143540 265032 143546
rect 264980 143482 265032 143488
rect 264428 132320 264480 132326
rect 264428 132262 264480 132268
rect 264518 131744 264574 131753
rect 264518 131679 264574 131688
rect 264336 118652 264388 118658
rect 264336 118594 264388 118600
rect 264244 117360 264296 117366
rect 264244 117302 264296 117308
rect 262864 46300 262916 46306
rect 262864 46242 262916 46248
rect 262220 28348 262272 28354
rect 262220 28290 262272 28296
rect 261484 22772 261536 22778
rect 261484 22714 261536 22720
rect 262232 16574 262260 28290
rect 260852 16546 261800 16574
rect 262232 16546 262536 16574
rect 259460 13184 259512 13190
rect 259460 13126 259512 13132
rect 258724 4820 258776 4826
rect 258724 4762 258776 4768
rect 259472 3602 259500 13126
rect 259460 3596 259512 3602
rect 259460 3538 259512 3544
rect 260656 3596 260708 3602
rect 260656 3538 260708 3544
rect 258262 3496 258318 3505
rect 258262 3431 258318 3440
rect 259458 3496 259514 3505
rect 259458 3431 259514 3440
rect 258276 480 258304 3431
rect 259472 480 259500 3431
rect 260668 480 260696 3538
rect 261772 480 261800 16546
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 264256 10402 264284 117302
rect 264532 99278 264560 131679
rect 265636 121378 265664 160142
rect 266464 155786 266492 185914
rect 266544 183048 266596 183054
rect 266544 182990 266596 182996
rect 266556 164218 266584 182990
rect 267004 172576 267056 172582
rect 267004 172518 267056 172524
rect 266544 164212 266596 164218
rect 266544 164154 266596 164160
rect 266452 155780 266504 155786
rect 266452 155722 266504 155728
rect 265716 135312 265768 135318
rect 265716 135254 265768 135260
rect 265624 121372 265676 121378
rect 265624 121314 265676 121320
rect 265624 117428 265676 117434
rect 265624 117370 265676 117376
rect 264520 99272 264572 99278
rect 264520 99214 264572 99220
rect 265636 26926 265664 117370
rect 265728 75274 265756 135254
rect 267016 133754 267044 172518
rect 267752 162790 267780 231066
rect 267924 188624 267976 188630
rect 267924 188566 267976 188572
rect 267832 180260 267884 180266
rect 267832 180202 267884 180208
rect 267740 162784 267792 162790
rect 267740 162726 267792 162732
rect 267096 154692 267148 154698
rect 267096 154634 267148 154640
rect 267004 133748 267056 133754
rect 267004 133690 267056 133696
rect 267004 121508 267056 121514
rect 267004 121450 267056 121456
rect 265716 75268 265768 75274
rect 265716 75210 265768 75216
rect 265624 26920 265676 26926
rect 265624 26862 265676 26868
rect 267016 19990 267044 121450
rect 267108 115938 267136 154634
rect 267844 144906 267872 180202
rect 267936 153134 267964 188566
rect 268384 171216 268436 171222
rect 268384 171158 268436 171164
rect 267924 153128 267976 153134
rect 267924 153070 267976 153076
rect 267832 144900 267884 144906
rect 267832 144842 267884 144848
rect 267188 139460 267240 139466
rect 267188 139402 267240 139408
rect 267096 115932 267148 115938
rect 267096 115874 267148 115880
rect 267200 101454 267228 139402
rect 268396 133822 268424 171158
rect 268476 156052 268528 156058
rect 268476 155994 268528 156000
rect 268384 133816 268436 133822
rect 268384 133758 268436 133764
rect 268488 117230 268516 155994
rect 268476 117224 268528 117230
rect 268476 117166 268528 117172
rect 268384 116000 268436 116006
rect 268384 115942 268436 115948
rect 267188 101448 267240 101454
rect 267188 101390 267240 101396
rect 267096 100972 267148 100978
rect 267096 100914 267148 100920
rect 267004 19984 267056 19990
rect 267004 19926 267056 19932
rect 267108 18698 267136 100914
rect 267096 18692 267148 18698
rect 267096 18634 267148 18640
rect 268396 15910 268424 115942
rect 269132 16574 269160 336126
rect 269776 291174 269804 349114
rect 269764 291168 269816 291174
rect 269764 291110 269816 291116
rect 270500 209160 270552 209166
rect 270500 209102 270552 209108
rect 269212 195424 269264 195430
rect 269212 195366 269264 195372
rect 269224 154494 269252 195366
rect 269764 173936 269816 173942
rect 269764 173878 269816 173884
rect 269212 154488 269264 154494
rect 269212 154430 269264 154436
rect 269776 136474 269804 173878
rect 270512 165578 270540 209102
rect 270684 199504 270736 199510
rect 270684 199446 270736 199452
rect 270592 184408 270644 184414
rect 270592 184350 270644 184356
rect 270500 165572 270552 165578
rect 270500 165514 270552 165520
rect 269856 164892 269908 164898
rect 269856 164834 269908 164840
rect 269764 136468 269816 136474
rect 269764 136410 269816 136416
rect 269868 131034 269896 164834
rect 270604 146198 270632 184350
rect 270696 161430 270724 199446
rect 271328 168496 271380 168502
rect 271328 168438 271380 168444
rect 271236 162988 271288 162994
rect 271236 162930 271288 162936
rect 270684 161424 270736 161430
rect 270684 161366 270736 161372
rect 270592 146192 270644 146198
rect 270592 146134 270644 146140
rect 269856 131028 269908 131034
rect 269856 130970 269908 130976
rect 269948 130416 270000 130422
rect 269948 130358 270000 130364
rect 269764 114572 269816 114578
rect 269764 114514 269816 114520
rect 269776 57254 269804 114514
rect 269960 100570 269988 130358
rect 271144 128376 271196 128382
rect 271144 128318 271196 128324
rect 269948 100564 270000 100570
rect 269948 100506 270000 100512
rect 269764 57248 269816 57254
rect 269764 57190 269816 57196
rect 271156 44946 271184 128318
rect 271248 124098 271276 162930
rect 271340 129674 271368 168438
rect 271328 129668 271380 129674
rect 271328 129610 271380 129616
rect 271236 124092 271288 124098
rect 271236 124034 271288 124040
rect 271236 120148 271288 120154
rect 271236 120090 271288 120096
rect 271248 72554 271276 120090
rect 271236 72548 271288 72554
rect 271236 72490 271288 72496
rect 271144 44940 271196 44946
rect 271144 44882 271196 44888
rect 270500 32428 270552 32434
rect 270500 32370 270552 32376
rect 270512 16574 270540 32370
rect 271892 16574 271920 370466
rect 278044 346452 278096 346458
rect 278044 346394 278096 346400
rect 277400 342916 277452 342922
rect 277400 342858 277452 342864
rect 273260 333260 273312 333266
rect 273260 333202 273312 333208
rect 272064 198144 272116 198150
rect 272064 198086 272116 198092
rect 271972 182980 272024 182986
rect 271972 182922 272024 182928
rect 271984 142118 272012 182922
rect 272076 157350 272104 198086
rect 272616 178084 272668 178090
rect 272616 178026 272668 178032
rect 272064 157344 272116 157350
rect 272064 157286 272116 157292
rect 271972 142112 272024 142118
rect 271972 142054 272024 142060
rect 272524 122868 272576 122874
rect 272524 122810 272576 122816
rect 272536 24138 272564 122810
rect 272628 97306 272656 178026
rect 272800 151904 272852 151910
rect 272800 151846 272852 151852
rect 272812 111722 272840 151846
rect 272800 111716 272852 111722
rect 272800 111658 272852 111664
rect 272708 110492 272760 110498
rect 272708 110434 272760 110440
rect 272616 97300 272668 97306
rect 272616 97242 272668 97248
rect 272720 53106 272748 110434
rect 272708 53100 272760 53106
rect 272708 53042 272760 53048
rect 272524 24132 272576 24138
rect 272524 24074 272576 24080
rect 269132 16546 270080 16574
rect 270512 16546 270816 16574
rect 271892 16546 272472 16574
rect 268384 15904 268436 15910
rect 268384 15846 268436 15852
rect 267740 13116 267792 13122
rect 267740 13058 267792 13064
rect 264244 10396 264296 10402
rect 264244 10338 264296 10344
rect 264150 3496 264206 3505
rect 264150 3431 264206 3440
rect 265346 3496 265402 3505
rect 265346 3431 265402 3440
rect 266542 3496 266598 3505
rect 266542 3431 266598 3440
rect 264164 480 264192 3431
rect 265360 480 265388 3431
rect 266556 480 266584 3431
rect 267752 480 267780 13058
rect 268842 3632 268898 3641
rect 268842 3567 268898 3576
rect 268856 480 268884 3567
rect 270052 480 270080 16546
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270788 354 270816 16546
rect 272444 480 272472 16546
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273272 354 273300 333202
rect 274640 308576 274692 308582
rect 274640 308518 274692 308524
rect 273902 293176 273958 293185
rect 273902 293111 273958 293120
rect 273916 259418 273944 293111
rect 273904 259412 273956 259418
rect 273904 259354 273956 259360
rect 273352 193928 273404 193934
rect 273352 193870 273404 193876
rect 273364 147558 273392 193870
rect 273536 181620 273588 181626
rect 273536 181562 273588 181568
rect 273444 180192 273496 180198
rect 273444 180134 273496 180140
rect 273352 147552 273404 147558
rect 273352 147494 273404 147500
rect 273456 137902 273484 180134
rect 273548 153202 273576 181562
rect 273536 153196 273588 153202
rect 273536 153138 273588 153144
rect 273996 150544 274048 150550
rect 273996 150486 274048 150492
rect 273444 137896 273496 137902
rect 273444 137838 273496 137844
rect 273904 132524 273956 132530
rect 273904 132466 273956 132472
rect 273916 72486 273944 132466
rect 274008 110362 274036 150486
rect 273996 110356 274048 110362
rect 273996 110298 274048 110304
rect 273996 100836 274048 100842
rect 273996 100778 274048 100784
rect 273904 72480 273956 72486
rect 273904 72422 273956 72428
rect 274008 43450 274036 100778
rect 273996 43444 274048 43450
rect 273996 43386 274048 43392
rect 274652 16574 274680 308518
rect 276112 292664 276164 292670
rect 276112 292606 276164 292612
rect 276020 291168 276072 291174
rect 276020 291110 276072 291116
rect 274824 198212 274876 198218
rect 274824 198154 274876 198160
rect 274732 185904 274784 185910
rect 274732 185846 274784 185852
rect 274744 139398 274772 185846
rect 274836 160070 274864 198154
rect 275376 169788 275428 169794
rect 275376 169730 275428 169736
rect 274824 160064 274876 160070
rect 274824 160006 274876 160012
rect 274732 139392 274784 139398
rect 274732 139334 274784 139340
rect 275388 131102 275416 169730
rect 275468 149728 275520 149734
rect 275468 149670 275520 149676
rect 275376 131096 275428 131102
rect 275376 131038 275428 131044
rect 275284 129804 275336 129810
rect 275284 129746 275336 129752
rect 275296 38010 275324 129746
rect 275480 114510 275508 149670
rect 275468 114504 275520 114510
rect 275468 114446 275520 114452
rect 275376 109064 275428 109070
rect 275376 109006 275428 109012
rect 275388 61470 275416 109006
rect 275376 61464 275428 61470
rect 275376 61406 275428 61412
rect 275284 38004 275336 38010
rect 275284 37946 275336 37952
rect 274652 16546 274864 16574
rect 274836 480 274864 16546
rect 276032 480 276060 291110
rect 276124 137970 276152 292606
rect 276204 187060 276256 187066
rect 276204 187002 276256 187008
rect 276216 158710 276244 187002
rect 276664 167068 276716 167074
rect 276664 167010 276716 167016
rect 276204 158704 276256 158710
rect 276204 158646 276256 158652
rect 276112 137964 276164 137970
rect 276112 137906 276164 137912
rect 276676 129742 276704 167010
rect 276756 142248 276808 142254
rect 276756 142190 276808 142196
rect 276664 129736 276716 129742
rect 276664 129678 276716 129684
rect 276664 113280 276716 113286
rect 276664 113222 276716 113228
rect 276676 60042 276704 113222
rect 276768 102134 276796 142190
rect 276756 102128 276808 102134
rect 276756 102070 276808 102076
rect 276664 60036 276716 60042
rect 276664 59978 276716 59984
rect 277412 16574 277440 342858
rect 277492 191344 277544 191350
rect 277492 191286 277544 191292
rect 277504 150414 277532 191286
rect 277492 150408 277544 150414
rect 277492 150350 277544 150356
rect 278056 61470 278084 346394
rect 278780 307080 278832 307086
rect 278780 307022 278832 307028
rect 278228 165708 278280 165714
rect 278228 165650 278280 165656
rect 278136 138100 278188 138106
rect 278136 138042 278188 138048
rect 278044 61464 278096 61470
rect 278044 61406 278096 61412
rect 277412 16546 278084 16574
rect 277122 3632 277178 3641
rect 277122 3567 277178 3576
rect 277136 480 277164 3567
rect 278056 3482 278084 16546
rect 278148 4894 278176 138042
rect 278240 128178 278268 165650
rect 278228 128172 278280 128178
rect 278228 128114 278280 128120
rect 278228 96756 278280 96762
rect 278228 96698 278280 96704
rect 278240 36582 278268 96698
rect 278228 36576 278280 36582
rect 278228 36518 278280 36524
rect 278792 16574 278820 307022
rect 279422 297392 279478 297401
rect 279422 297327 279478 297336
rect 278872 207664 278924 207670
rect 278872 207606 278924 207612
rect 278884 148986 278912 207606
rect 278872 148980 278924 148986
rect 278872 148922 278924 148928
rect 278792 16546 279096 16574
rect 278136 4888 278188 4894
rect 278136 4830 278188 4836
rect 278056 3454 278360 3482
rect 278332 480 278360 3454
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 279436 3466 279464 297327
rect 280160 214668 280212 214674
rect 280160 214610 280212 214616
rect 280172 146266 280200 214610
rect 280252 192636 280304 192642
rect 280252 192578 280304 192584
rect 280264 149054 280292 192578
rect 280252 149048 280304 149054
rect 280252 148990 280304 148996
rect 280160 146260 280212 146266
rect 280160 146202 280212 146208
rect 279608 144968 279660 144974
rect 279608 144910 279660 144916
rect 279620 104174 279648 144910
rect 279608 104168 279660 104174
rect 279608 104110 279660 104116
rect 279516 103556 279568 103562
rect 279516 103498 279568 103504
rect 279528 39438 279556 103498
rect 280816 78062 280844 382570
rect 282920 363656 282972 363662
rect 282920 363598 282972 363604
rect 281540 329112 281592 329118
rect 281540 329054 281592 329060
rect 281080 167136 281132 167142
rect 281080 167078 281132 167084
rect 280896 128444 280948 128450
rect 280896 128386 280948 128392
rect 280804 78056 280856 78062
rect 280804 77998 280856 78004
rect 280908 40798 280936 128386
rect 281092 128246 281120 167078
rect 281080 128240 281132 128246
rect 281080 128182 281132 128188
rect 280988 127016 281040 127022
rect 280988 126958 281040 126964
rect 281000 42158 281028 126958
rect 280988 42152 281040 42158
rect 280988 42094 281040 42100
rect 280896 40792 280948 40798
rect 280896 40734 280948 40740
rect 279516 39432 279568 39438
rect 279516 39374 279568 39380
rect 280160 21412 280212 21418
rect 280160 21354 280212 21360
rect 280172 16574 280200 21354
rect 280172 16546 280752 16574
rect 279424 3460 279476 3466
rect 279424 3402 279476 3408
rect 280724 480 280752 16546
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281552 354 281580 329054
rect 281632 205012 281684 205018
rect 281632 204954 281684 204960
rect 281644 151774 281672 204954
rect 281724 189916 281776 189922
rect 281724 189858 281776 189864
rect 281632 151768 281684 151774
rect 281632 151710 281684 151716
rect 281736 140758 281764 189858
rect 282460 155236 282512 155242
rect 282460 155178 282512 155184
rect 281724 140752 281776 140758
rect 281724 140694 281776 140700
rect 282276 139528 282328 139534
rect 282276 139470 282328 139476
rect 282184 127084 282236 127090
rect 282184 127026 282236 127032
rect 282196 6186 282224 127026
rect 282288 51814 282316 139470
rect 282472 117298 282500 155178
rect 282460 117292 282512 117298
rect 282460 117234 282512 117240
rect 282368 116068 282420 116074
rect 282368 116010 282420 116016
rect 282380 61402 282408 116010
rect 282368 61396 282420 61402
rect 282368 61338 282420 61344
rect 282276 51808 282328 51814
rect 282276 51750 282328 51756
rect 282932 16574 282960 363598
rect 284300 338768 284352 338774
rect 284300 338710 284352 338716
rect 283748 167204 283800 167210
rect 283748 167146 283800 167152
rect 283564 131164 283616 131170
rect 283564 131106 283616 131112
rect 283576 33794 283604 131106
rect 283760 128314 283788 167146
rect 283748 128308 283800 128314
rect 283748 128250 283800 128256
rect 283656 127152 283708 127158
rect 283656 127094 283708 127100
rect 283668 39370 283696 127094
rect 283656 39364 283708 39370
rect 283656 39306 283708 39312
rect 283564 33788 283616 33794
rect 283564 33730 283616 33736
rect 282932 16546 283144 16574
rect 282184 6180 282236 6186
rect 282184 6122 282236 6128
rect 283116 480 283144 16546
rect 284312 480 284340 338710
rect 307024 337408 307076 337414
rect 307024 337350 307076 337356
rect 293960 330540 294012 330546
rect 293960 330482 294012 330488
rect 284392 323672 284444 323678
rect 284392 323614 284444 323620
rect 284404 16574 284432 323614
rect 287060 322312 287112 322318
rect 287060 322254 287112 322260
rect 286324 236700 286376 236706
rect 286324 236642 286376 236648
rect 285036 135380 285088 135386
rect 285036 135322 285088 135328
rect 284944 113348 284996 113354
rect 284944 113290 284996 113296
rect 284956 49026 284984 113290
rect 285048 73914 285076 135322
rect 286336 96558 286364 236642
rect 286416 169856 286468 169862
rect 286416 169798 286468 169804
rect 286428 132394 286456 169798
rect 286692 134564 286744 134570
rect 286692 134506 286744 134512
rect 286416 132388 286468 132394
rect 286416 132330 286468 132336
rect 286508 131232 286560 131238
rect 286508 131174 286560 131180
rect 286416 120216 286468 120222
rect 286416 120158 286468 120164
rect 286324 96552 286376 96558
rect 286324 96494 286376 96500
rect 285036 73908 285088 73914
rect 285036 73850 285088 73856
rect 284944 49020 284996 49026
rect 284944 48962 284996 48968
rect 284404 16546 284984 16574
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 354 284984 16546
rect 286428 11762 286456 120158
rect 286520 65550 286548 131174
rect 286704 99210 286732 134506
rect 286692 99204 286744 99210
rect 286692 99146 286744 99152
rect 286600 98116 286652 98122
rect 286600 98058 286652 98064
rect 286508 65544 286560 65550
rect 286508 65486 286560 65492
rect 286612 37942 286640 98058
rect 286600 37936 286652 37942
rect 286600 37878 286652 37884
rect 287072 16574 287100 322254
rect 287704 312656 287756 312662
rect 287704 312598 287756 312604
rect 287072 16546 287376 16574
rect 286416 11756 286468 11762
rect 286416 11698 286468 11704
rect 286598 3496 286654 3505
rect 286598 3431 286654 3440
rect 286612 480 286640 3431
rect 285374 354 285486 480
rect 284956 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 287716 3534 287744 312598
rect 291200 309800 291252 309806
rect 291200 309742 291252 309748
rect 289176 174004 289228 174010
rect 289176 173946 289228 173952
rect 289084 172644 289136 172650
rect 289084 172586 289136 172592
rect 287980 164280 288032 164286
rect 287980 164222 288032 164228
rect 287796 132592 287848 132598
rect 287796 132534 287848 132540
rect 287808 31074 287836 132534
rect 287992 125526 288020 164222
rect 289096 135182 289124 172586
rect 289188 136542 289216 173946
rect 290464 168564 290516 168570
rect 290464 168506 290516 168512
rect 290476 140078 290504 168506
rect 290740 144288 290792 144294
rect 290740 144230 290792 144236
rect 290464 140072 290516 140078
rect 290464 140014 290516 140020
rect 289176 136536 289228 136542
rect 289176 136478 289228 136484
rect 289268 135448 289320 135454
rect 289268 135390 289320 135396
rect 289084 135176 289136 135182
rect 289084 135118 289136 135124
rect 287980 125520 288032 125526
rect 287980 125462 288032 125468
rect 287888 124296 287940 124302
rect 287888 124238 287940 124244
rect 287900 35290 287928 124238
rect 289084 122936 289136 122942
rect 289084 122878 289136 122884
rect 287888 35284 287940 35290
rect 287888 35226 287940 35232
rect 287796 31068 287848 31074
rect 287796 31010 287848 31016
rect 289096 7614 289124 122878
rect 289176 102332 289228 102338
rect 289176 102274 289228 102280
rect 289188 10334 289216 102274
rect 289280 43518 289308 135390
rect 290648 129872 290700 129878
rect 290648 129814 290700 129820
rect 290556 128512 290608 128518
rect 290556 128454 290608 128460
rect 289360 125724 289412 125730
rect 289360 125666 289412 125672
rect 289372 66910 289400 125666
rect 290464 103624 290516 103630
rect 290464 103566 290516 103572
rect 289360 66904 289412 66910
rect 289360 66846 289412 66852
rect 289268 43512 289320 43518
rect 289268 43454 289320 43460
rect 290476 14482 290504 103566
rect 290568 47666 290596 128454
rect 290660 58682 290688 129814
rect 290752 104854 290780 144230
rect 290740 104848 290792 104854
rect 290740 104790 290792 104796
rect 290648 58676 290700 58682
rect 290648 58618 290700 58624
rect 290556 47660 290608 47666
rect 290556 47602 290608 47608
rect 291212 16574 291240 309742
rect 291936 174072 291988 174078
rect 291936 174014 291988 174020
rect 291844 160268 291896 160274
rect 291844 160210 291896 160216
rect 291856 121446 291884 160210
rect 291948 136610 291976 174014
rect 293408 157548 293460 157554
rect 293408 157490 293460 157496
rect 292028 136740 292080 136746
rect 292028 136682 292080 136688
rect 291936 136604 291988 136610
rect 291936 136546 291988 136552
rect 291844 121440 291896 121446
rect 291844 121382 291896 121388
rect 291844 118788 291896 118794
rect 291844 118730 291896 118736
rect 291856 22846 291884 118730
rect 291936 96824 291988 96830
rect 291936 96766 291988 96772
rect 291844 22840 291896 22846
rect 291844 22782 291896 22788
rect 291212 16546 291424 16574
rect 290464 14476 290516 14482
rect 290464 14418 290516 14424
rect 289176 10328 289228 10334
rect 289176 10270 289228 10276
rect 289084 7608 289136 7614
rect 289084 7550 289136 7556
rect 290186 3632 290242 3641
rect 290186 3567 290242 3576
rect 287704 3528 287756 3534
rect 287704 3470 287756 3476
rect 288990 3496 289046 3505
rect 288990 3431 289046 3440
rect 289004 480 289032 3431
rect 290200 480 290228 3567
rect 291396 480 291424 16546
rect 291948 2106 291976 96766
rect 292040 69766 292068 136682
rect 293224 133952 293276 133958
rect 293224 133894 293276 133900
rect 292028 69760 292080 69766
rect 292028 69702 292080 69708
rect 293236 50454 293264 133894
rect 293316 121576 293368 121582
rect 293316 121518 293368 121524
rect 293224 50448 293276 50454
rect 293224 50390 293276 50396
rect 293328 46238 293356 121518
rect 293420 119406 293448 157490
rect 293408 119400 293460 119406
rect 293408 119342 293460 119348
rect 293408 100904 293460 100910
rect 293408 100846 293460 100852
rect 293316 46232 293368 46238
rect 293316 46174 293368 46180
rect 293420 44878 293448 100846
rect 293408 44872 293460 44878
rect 293408 44814 293460 44820
rect 292580 24200 292632 24206
rect 292580 24142 292632 24148
rect 292592 16574 292620 24142
rect 293972 16574 294000 330482
rect 295984 310548 296036 310554
rect 295984 310490 296036 310496
rect 295996 180169 296024 310490
rect 298100 308508 298152 308514
rect 298100 308450 298152 308456
rect 296076 220108 296128 220114
rect 296076 220050 296128 220056
rect 295982 180160 296038 180169
rect 295982 180095 296038 180104
rect 296088 175817 296116 220050
rect 296074 175808 296130 175817
rect 296074 175743 296130 175752
rect 295984 172712 296036 172718
rect 295984 172654 296036 172660
rect 294880 141432 294932 141438
rect 294880 141374 294932 141380
rect 294604 138168 294656 138174
rect 294604 138110 294656 138116
rect 294616 68474 294644 138110
rect 294696 114640 294748 114646
rect 294696 114582 294748 114588
rect 294604 68468 294656 68474
rect 294604 68410 294656 68416
rect 294708 55894 294736 114582
rect 294892 100638 294920 141374
rect 295996 135250 296024 172654
rect 296076 171284 296128 171290
rect 296076 171226 296128 171232
rect 295984 135244 296036 135250
rect 295984 135186 296036 135192
rect 296088 133890 296116 171226
rect 297456 161628 297508 161634
rect 297456 161570 297508 161576
rect 296168 151972 296220 151978
rect 296168 151914 296220 151920
rect 296076 133884 296128 133890
rect 296076 133826 296128 133832
rect 295984 132660 296036 132666
rect 295984 132602 296036 132608
rect 294880 100632 294932 100638
rect 294880 100574 294932 100580
rect 294788 99408 294840 99414
rect 294788 99350 294840 99356
rect 294696 55888 294748 55894
rect 294696 55830 294748 55836
rect 294800 47598 294828 99350
rect 294788 47592 294840 47598
rect 294788 47534 294840 47540
rect 295996 17270 296024 132602
rect 296076 120284 296128 120290
rect 296076 120226 296128 120232
rect 296088 32502 296116 120226
rect 296180 111790 296208 151914
rect 297468 122806 297496 161570
rect 297640 153332 297692 153338
rect 297640 153274 297692 153280
rect 297456 122800 297508 122806
rect 297456 122742 297508 122748
rect 297364 121644 297416 121650
rect 297364 121586 297416 121592
rect 296352 116612 296404 116618
rect 296352 116554 296404 116560
rect 296168 111784 296220 111790
rect 296168 111726 296220 111732
rect 296260 110560 296312 110566
rect 296260 110502 296312 110508
rect 296168 99476 296220 99482
rect 296168 99418 296220 99424
rect 296180 40730 296208 99418
rect 296272 55962 296300 110502
rect 296364 100706 296392 116554
rect 296352 100700 296404 100706
rect 296352 100642 296404 100648
rect 296260 55956 296312 55962
rect 296260 55898 296312 55904
rect 296168 40724 296220 40730
rect 296168 40666 296220 40672
rect 296718 33824 296774 33833
rect 296718 33759 296774 33768
rect 296076 32496 296128 32502
rect 296076 32438 296128 32444
rect 295984 17264 296036 17270
rect 295984 17206 296036 17212
rect 296732 16574 296760 33759
rect 297376 25634 297404 121586
rect 297652 115258 297680 153274
rect 297732 149184 297784 149190
rect 297732 149126 297784 149132
rect 297640 115252 297692 115258
rect 297640 115194 297692 115200
rect 297548 114708 297600 114714
rect 297548 114650 297600 114656
rect 297456 111852 297508 111858
rect 297456 111794 297508 111800
rect 297468 26994 297496 111794
rect 297560 54534 297588 114650
rect 297744 108934 297772 149126
rect 297732 108928 297784 108934
rect 297732 108870 297784 108876
rect 297640 107908 297692 107914
rect 297640 107850 297692 107856
rect 297652 62830 297680 107850
rect 297640 62824 297692 62830
rect 297640 62766 297692 62772
rect 297548 54528 297600 54534
rect 297548 54470 297600 54476
rect 297456 26988 297508 26994
rect 297456 26930 297508 26936
rect 297364 25628 297416 25634
rect 297364 25570 297416 25576
rect 292592 16546 293264 16574
rect 293972 16546 294920 16574
rect 296732 16546 297312 16574
rect 292580 6316 292632 6322
rect 292580 6258 292632 6264
rect 291936 2100 291988 2106
rect 291936 2042 291988 2048
rect 292592 480 292620 6258
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 294892 480 294920 16546
rect 295616 16040 295668 16046
rect 295616 15982 295668 15988
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 295628 354 295656 15982
rect 297284 480 297312 16546
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298112 354 298140 308450
rect 300124 306400 300176 306406
rect 300124 306342 300176 306348
rect 300136 180198 300164 306342
rect 300216 217320 300268 217326
rect 300216 217262 300268 217268
rect 300124 180192 300176 180198
rect 300124 180134 300176 180140
rect 300228 180033 300256 217262
rect 300214 180024 300270 180033
rect 300214 179959 300270 179968
rect 307036 177410 307064 337350
rect 308404 322244 308456 322250
rect 308404 322186 308456 322192
rect 307116 260908 307168 260914
rect 307116 260850 307168 260856
rect 307128 182986 307156 260850
rect 307116 182980 307168 182986
rect 307116 182922 307168 182928
rect 307024 177404 307076 177410
rect 307024 177346 307076 177352
rect 307482 174856 307538 174865
rect 307482 174791 307538 174800
rect 307496 174010 307524 174791
rect 307574 174448 307630 174457
rect 307574 174383 307630 174392
rect 307484 174004 307536 174010
rect 307484 173946 307536 173952
rect 307588 173942 307616 174383
rect 307668 174072 307720 174078
rect 307666 174040 307668 174049
rect 307720 174040 307722 174049
rect 307666 173975 307722 173984
rect 307576 173936 307628 173942
rect 307576 173878 307628 173884
rect 307574 173632 307630 173641
rect 307574 173567 307630 173576
rect 307482 173224 307538 173233
rect 307482 173159 307538 173168
rect 307496 172718 307524 173159
rect 307484 172712 307536 172718
rect 307484 172654 307536 172660
rect 307588 172650 307616 173567
rect 307666 172680 307722 172689
rect 307576 172644 307628 172650
rect 307666 172615 307722 172624
rect 307576 172586 307628 172592
rect 307680 172582 307708 172615
rect 307668 172576 307720 172582
rect 307668 172518 307720 172524
rect 306562 172272 306618 172281
rect 306562 172207 306618 172216
rect 306576 171290 306604 172207
rect 307574 171864 307630 171873
rect 307574 171799 307630 171808
rect 306564 171284 306616 171290
rect 306564 171226 306616 171232
rect 307588 171222 307616 171799
rect 307666 171456 307722 171465
rect 307666 171391 307722 171400
rect 307576 171216 307628 171222
rect 307576 171158 307628 171164
rect 307680 171154 307708 171391
rect 307668 171148 307720 171154
rect 307668 171090 307720 171096
rect 307298 171048 307354 171057
rect 307298 170983 307354 170992
rect 300124 169924 300176 169930
rect 300124 169866 300176 169872
rect 298836 159384 298888 159390
rect 298836 159326 298888 159332
rect 298848 125594 298876 159326
rect 300136 132462 300164 169866
rect 307312 169862 307340 170983
rect 307666 170640 307722 170649
rect 307666 170575 307722 170584
rect 307482 170232 307538 170241
rect 307482 170167 307538 170176
rect 307300 169856 307352 169862
rect 307300 169798 307352 169804
rect 307390 169824 307446 169833
rect 307496 169794 307524 170167
rect 307680 169930 307708 170575
rect 307668 169924 307720 169930
rect 307668 169866 307720 169872
rect 307390 169759 307446 169768
rect 307484 169788 307536 169794
rect 307116 168564 307168 168570
rect 307116 168506 307168 168512
rect 307128 168473 307156 168506
rect 307114 168464 307170 168473
rect 307114 168399 307170 168408
rect 307298 168056 307354 168065
rect 307298 167991 307354 168000
rect 307312 167074 307340 167991
rect 307300 167068 307352 167074
rect 307300 167010 307352 167016
rect 307114 166424 307170 166433
rect 307114 166359 307170 166368
rect 307128 165782 307156 166359
rect 302884 165776 302936 165782
rect 302884 165718 302936 165724
rect 307116 165776 307168 165782
rect 307116 165718 307168 165724
rect 301504 163056 301556 163062
rect 301504 162998 301556 163004
rect 300768 156120 300820 156126
rect 300768 156062 300820 156068
rect 300780 153882 300808 156062
rect 300768 153876 300820 153882
rect 300768 153818 300820 153824
rect 300400 153400 300452 153406
rect 300400 153342 300452 153348
rect 300308 150612 300360 150618
rect 300308 150554 300360 150560
rect 300216 135516 300268 135522
rect 300216 135458 300268 135464
rect 300124 132456 300176 132462
rect 300124 132398 300176 132404
rect 298836 125588 298888 125594
rect 298836 125530 298888 125536
rect 298744 124364 298796 124370
rect 298744 124306 298796 124312
rect 298756 9042 298784 124306
rect 300124 117564 300176 117570
rect 300124 117506 300176 117512
rect 298836 117496 298888 117502
rect 298836 117438 298888 117444
rect 298848 18630 298876 117438
rect 298928 109132 298980 109138
rect 298928 109074 298980 109080
rect 298940 58750 298968 109074
rect 298928 58744 298980 58750
rect 298928 58686 298980 58692
rect 300136 21486 300164 117506
rect 300228 76566 300256 135458
rect 300320 110430 300348 150554
rect 300412 113150 300440 153342
rect 301516 124166 301544 162998
rect 301780 146668 301832 146674
rect 301780 146610 301832 146616
rect 301504 124160 301556 124166
rect 301504 124102 301556 124108
rect 301688 123004 301740 123010
rect 301688 122946 301740 122952
rect 300400 113144 300452 113150
rect 300400 113086 300452 113092
rect 301504 111988 301556 111994
rect 301504 111930 301556 111936
rect 300308 110424 300360 110430
rect 300308 110366 300360 110372
rect 300400 107772 300452 107778
rect 300400 107714 300452 107720
rect 300308 99544 300360 99550
rect 300308 99486 300360 99492
rect 300216 76560 300268 76566
rect 300216 76502 300268 76508
rect 300320 51746 300348 99486
rect 300412 66978 300440 107714
rect 300400 66972 300452 66978
rect 300400 66914 300452 66920
rect 300308 51740 300360 51746
rect 300308 51682 300360 51688
rect 301516 28286 301544 111930
rect 301596 109200 301648 109206
rect 301596 109142 301648 109148
rect 301608 57322 301636 109142
rect 301700 71126 301728 122946
rect 301792 109002 301820 146610
rect 302896 126954 302924 165718
rect 307022 165472 307078 165481
rect 307022 165407 307078 165416
rect 305736 164348 305788 164354
rect 305736 164290 305788 164296
rect 305642 147792 305698 147801
rect 305642 147727 305698 147736
rect 304356 147688 304408 147694
rect 304356 147630 304408 147636
rect 303068 145036 303120 145042
rect 303068 144978 303120 144984
rect 302884 126948 302936 126954
rect 302884 126890 302936 126896
rect 302884 124432 302936 124438
rect 302884 124374 302936 124380
rect 301780 108996 301832 109002
rect 301780 108938 301832 108944
rect 301780 106412 301832 106418
rect 301780 106354 301832 106360
rect 301688 71120 301740 71126
rect 301688 71062 301740 71068
rect 301792 68406 301820 106354
rect 301780 68400 301832 68406
rect 301780 68342 301832 68348
rect 301596 57316 301648 57322
rect 301596 57258 301648 57264
rect 301504 28280 301556 28286
rect 301504 28222 301556 28228
rect 300124 21480 300176 21486
rect 300124 21422 300176 21428
rect 298836 18624 298888 18630
rect 298836 18566 298888 18572
rect 302896 17338 302924 124374
rect 303080 112470 303108 144978
rect 304264 118856 304316 118862
rect 304264 118798 304316 118804
rect 303068 112464 303120 112470
rect 303068 112406 303120 112412
rect 302976 111920 303028 111926
rect 302976 111862 303028 111868
rect 302988 49094 303016 111862
rect 303068 107704 303120 107710
rect 303068 107646 303120 107652
rect 303080 64190 303108 107646
rect 303160 104916 303212 104922
rect 303160 104858 303212 104864
rect 303172 75206 303200 104858
rect 303160 75200 303212 75206
rect 303160 75142 303212 75148
rect 303068 64184 303120 64190
rect 303068 64126 303120 64132
rect 302976 49088 303028 49094
rect 302976 49030 303028 49036
rect 302884 17332 302936 17338
rect 302884 17274 302936 17280
rect 299478 14512 299534 14521
rect 299478 14447 299534 14456
rect 298744 9036 298796 9042
rect 298744 8978 298796 8984
rect 299492 3602 299520 14447
rect 299480 3596 299532 3602
rect 299480 3538 299532 3544
rect 300768 3596 300820 3602
rect 300768 3538 300820 3544
rect 299662 3360 299718 3369
rect 299662 3295 299718 3304
rect 299676 480 299704 3295
rect 300780 480 300808 3538
rect 301962 3496 302018 3505
rect 301962 3431 302018 3440
rect 303158 3496 303214 3505
rect 303158 3431 303214 3440
rect 301976 480 302004 3431
rect 303172 480 303200 3431
rect 304276 2174 304304 118798
rect 304368 107574 304396 147630
rect 304540 143676 304592 143682
rect 304540 143618 304592 143624
rect 304448 110628 304500 110634
rect 304448 110570 304500 110576
rect 304356 107568 304408 107574
rect 304356 107510 304408 107516
rect 304356 103692 304408 103698
rect 304356 103634 304408 103640
rect 304368 25566 304396 103634
rect 304460 54602 304488 110570
rect 304552 105602 304580 143618
rect 305656 107642 305684 147727
rect 305748 126274 305776 164290
rect 306746 163432 306802 163441
rect 306746 163367 306802 163376
rect 306760 162994 306788 163367
rect 306748 162988 306800 162994
rect 306748 162930 306800 162936
rect 306562 161256 306618 161265
rect 306562 161191 306618 161200
rect 306576 160206 306604 161191
rect 306564 160200 306616 160206
rect 306564 160142 306616 160148
rect 306930 158672 306986 158681
rect 306930 158607 306986 158616
rect 306944 157486 306972 158607
rect 306932 157480 306984 157486
rect 306932 157422 306984 157428
rect 306562 155680 306618 155689
rect 306562 155615 306618 155624
rect 306576 154698 306604 155615
rect 306564 154692 306616 154698
rect 306564 154634 306616 154640
rect 306562 154456 306618 154465
rect 306562 154391 306618 154400
rect 306576 153270 306604 154391
rect 306564 153264 306616 153270
rect 306564 153206 306616 153212
rect 306654 153232 306710 153241
rect 306654 153167 306710 153176
rect 306562 152688 306618 152697
rect 306562 152623 306618 152632
rect 306576 151978 306604 152623
rect 306564 151972 306616 151978
rect 306564 151914 306616 151920
rect 306562 149832 306618 149841
rect 306562 149767 306618 149776
rect 306576 149122 306604 149767
rect 306564 149116 306616 149122
rect 306564 149058 306616 149064
rect 306668 148374 306696 153167
rect 306656 148368 306708 148374
rect 306656 148310 306708 148316
rect 306930 146840 306986 146849
rect 306930 146775 306986 146784
rect 306746 146432 306802 146441
rect 306746 146367 306802 146376
rect 306562 144664 306618 144673
rect 306562 144599 306618 144608
rect 306576 143614 306604 144599
rect 306654 143848 306710 143857
rect 306654 143783 306710 143792
rect 306564 143608 306616 143614
rect 306564 143550 306616 143556
rect 306470 142488 306526 142497
rect 306470 142423 306526 142432
rect 306484 141438 306512 142423
rect 306668 141545 306696 143783
rect 306760 142769 306788 146367
rect 306944 146334 306972 146775
rect 306932 146328 306984 146334
rect 306932 146270 306984 146276
rect 306746 142760 306802 142769
rect 306746 142695 306802 142704
rect 306654 141536 306710 141545
rect 306654 141471 306710 141480
rect 306472 141432 306524 141438
rect 306472 141374 306524 141380
rect 307036 137290 307064 165407
rect 307114 165064 307170 165073
rect 307114 164999 307170 165008
rect 307128 164354 307156 164999
rect 307404 164898 307432 169759
rect 307484 169730 307536 169736
rect 307574 169280 307630 169289
rect 307574 169215 307630 169224
rect 307588 168434 307616 169215
rect 307666 168872 307722 168881
rect 307666 168807 307722 168816
rect 307680 168502 307708 168807
rect 307668 168496 307720 168502
rect 307668 168438 307720 168444
rect 307576 168428 307628 168434
rect 307576 168370 307628 168376
rect 307482 167648 307538 167657
rect 307482 167583 307538 167592
rect 307496 167210 307524 167583
rect 307666 167240 307722 167249
rect 307484 167204 307536 167210
rect 307666 167175 307722 167184
rect 307484 167146 307536 167152
rect 307680 167142 307708 167175
rect 307668 167136 307720 167142
rect 307668 167078 307720 167084
rect 307574 166832 307630 166841
rect 307574 166767 307630 166776
rect 307588 165714 307616 166767
rect 307666 165880 307722 165889
rect 307666 165815 307722 165824
rect 307576 165708 307628 165714
rect 307576 165650 307628 165656
rect 307680 165646 307708 165815
rect 307668 165640 307720 165646
rect 307668 165582 307720 165588
rect 307392 164892 307444 164898
rect 307392 164834 307444 164840
rect 307206 164656 307262 164665
rect 307206 164591 307262 164600
rect 307116 164348 307168 164354
rect 307116 164290 307168 164296
rect 307114 159624 307170 159633
rect 307114 159559 307170 159568
rect 307128 145586 307156 159559
rect 307220 159390 307248 164591
rect 307668 164280 307720 164286
rect 307666 164248 307668 164257
rect 307720 164248 307722 164257
rect 307666 164183 307722 164192
rect 307574 163840 307630 163849
rect 307574 163775 307630 163784
rect 307588 163062 307616 163775
rect 307576 163056 307628 163062
rect 307576 162998 307628 163004
rect 307666 163024 307722 163033
rect 307666 162959 307722 162968
rect 307680 162926 307708 162959
rect 307668 162920 307720 162926
rect 307668 162862 307720 162868
rect 307482 162480 307538 162489
rect 307482 162415 307538 162424
rect 307496 161634 307524 162415
rect 307574 162072 307630 162081
rect 307574 162007 307630 162016
rect 307484 161628 307536 161634
rect 307484 161570 307536 161576
rect 307588 161566 307616 162007
rect 307666 161664 307722 161673
rect 307666 161599 307722 161608
rect 307576 161560 307628 161566
rect 307576 161502 307628 161508
rect 307680 161498 307708 161599
rect 307668 161492 307720 161498
rect 307668 161434 307720 161440
rect 307666 160848 307722 160857
rect 307666 160783 307722 160792
rect 307574 160440 307630 160449
rect 307574 160375 307630 160384
rect 307588 160138 307616 160375
rect 307680 160274 307708 160783
rect 307668 160268 307720 160274
rect 307668 160210 307720 160216
rect 307576 160132 307628 160138
rect 307576 160074 307628 160080
rect 307574 160032 307630 160041
rect 307574 159967 307630 159976
rect 307208 159384 307260 159390
rect 307208 159326 307260 159332
rect 307588 158846 307616 159967
rect 307666 159080 307722 159089
rect 307666 159015 307722 159024
rect 307576 158840 307628 158846
rect 307576 158782 307628 158788
rect 307680 158778 307708 159015
rect 307668 158772 307720 158778
rect 307668 158714 307720 158720
rect 307574 158264 307630 158273
rect 307574 158199 307630 158208
rect 307390 157448 307446 157457
rect 307588 157418 307616 158199
rect 307666 157856 307722 157865
rect 307666 157791 307722 157800
rect 307680 157554 307708 157791
rect 307668 157548 307720 157554
rect 307668 157490 307720 157496
rect 307390 157383 307446 157392
rect 307576 157412 307628 157418
rect 307404 155242 307432 157383
rect 307576 157354 307628 157360
rect 307482 157040 307538 157049
rect 307482 156975 307538 156984
rect 307496 156058 307524 156975
rect 307574 156632 307630 156641
rect 307574 156567 307630 156576
rect 307484 156052 307536 156058
rect 307484 155994 307536 156000
rect 307588 155990 307616 156567
rect 307666 156224 307722 156233
rect 307666 156159 307722 156168
rect 307680 156126 307708 156159
rect 307668 156120 307720 156126
rect 307668 156062 307720 156068
rect 307576 155984 307628 155990
rect 307576 155926 307628 155932
rect 307666 155272 307722 155281
rect 307392 155236 307444 155242
rect 307666 155207 307722 155216
rect 307392 155178 307444 155184
rect 307206 154864 307262 154873
rect 307206 154799 307262 154808
rect 307220 149734 307248 154799
rect 307680 154630 307708 155207
rect 307668 154624 307720 154630
rect 307668 154566 307720 154572
rect 307574 154048 307630 154057
rect 307574 153983 307630 153992
rect 307588 153406 307616 153983
rect 307666 153640 307722 153649
rect 307666 153575 307722 153584
rect 307576 153400 307628 153406
rect 307576 153342 307628 153348
rect 307680 153338 307708 153575
rect 307668 153332 307720 153338
rect 307668 153274 307720 153280
rect 307482 152280 307538 152289
rect 307482 152215 307538 152224
rect 307496 151842 307524 152215
rect 307668 151904 307720 151910
rect 307666 151872 307668 151881
rect 307720 151872 307722 151881
rect 307484 151836 307536 151842
rect 307666 151807 307722 151816
rect 307484 151778 307536 151784
rect 307482 151464 307538 151473
rect 307482 151399 307538 151408
rect 307496 150550 307524 151399
rect 307666 151056 307722 151065
rect 307666 150991 307722 151000
rect 307574 150648 307630 150657
rect 307680 150618 307708 150991
rect 307574 150583 307630 150592
rect 307668 150612 307720 150618
rect 307484 150544 307536 150550
rect 307484 150486 307536 150492
rect 307588 150482 307616 150583
rect 307668 150554 307720 150560
rect 307576 150476 307628 150482
rect 307576 150418 307628 150424
rect 307482 150240 307538 150249
rect 307482 150175 307538 150184
rect 307208 149728 307260 149734
rect 307208 149670 307260 149676
rect 307496 149190 307524 150175
rect 307574 149288 307630 149297
rect 307574 149223 307630 149232
rect 307484 149184 307536 149190
rect 307484 149126 307536 149132
rect 307298 148880 307354 148889
rect 307298 148815 307354 148824
rect 307312 147694 307340 148815
rect 307300 147688 307352 147694
rect 307300 147630 307352 147636
rect 307390 147656 307446 147665
rect 307390 147591 307446 147600
rect 307298 147248 307354 147257
rect 307298 147183 307354 147192
rect 307312 146402 307340 147183
rect 307300 146396 307352 146402
rect 307300 146338 307352 146344
rect 307116 145580 307168 145586
rect 307116 145522 307168 145528
rect 307404 144226 307432 147591
rect 307588 146674 307616 149223
rect 307666 148472 307722 148481
rect 307666 148407 307722 148416
rect 307680 147830 307708 148407
rect 307668 147824 307720 147830
rect 307668 147766 307720 147772
rect 307576 146668 307628 146674
rect 307576 146610 307628 146616
rect 307574 145888 307630 145897
rect 307574 145823 307630 145832
rect 307482 145480 307538 145489
rect 307482 145415 307538 145424
rect 307496 145042 307524 145415
rect 307484 145036 307536 145042
rect 307484 144978 307536 144984
rect 307588 144294 307616 145823
rect 307666 145072 307722 145081
rect 307666 145007 307722 145016
rect 307680 144974 307708 145007
rect 307668 144968 307720 144974
rect 307668 144910 307720 144916
rect 307576 144288 307628 144294
rect 307576 144230 307628 144236
rect 307666 144256 307722 144265
rect 307392 144220 307444 144226
rect 307666 144191 307722 144200
rect 307392 144162 307444 144168
rect 307680 143682 307708 144191
rect 307668 143676 307720 143682
rect 307668 143618 307720 143624
rect 307574 143440 307630 143449
rect 307574 143375 307630 143384
rect 307588 142186 307616 143375
rect 307666 143032 307722 143041
rect 307666 142967 307722 142976
rect 307680 142254 307708 142967
rect 307668 142248 307720 142254
rect 307668 142190 307720 142196
rect 307576 142180 307628 142186
rect 307576 142122 307628 142128
rect 307206 142080 307262 142089
rect 307206 142015 307262 142024
rect 307114 141672 307170 141681
rect 307114 141607 307170 141616
rect 307024 137284 307076 137290
rect 307024 137226 307076 137232
rect 306746 135688 306802 135697
rect 306746 135623 306802 135632
rect 306760 135522 306788 135623
rect 306748 135516 306800 135522
rect 306748 135458 306800 135464
rect 306562 133648 306618 133657
rect 306562 133583 306618 133592
rect 306576 132666 306604 133583
rect 307128 133362 307156 141607
rect 307220 137170 307248 142015
rect 307390 140856 307446 140865
rect 307390 140791 307446 140800
rect 307298 139632 307354 139641
rect 307298 139567 307354 139576
rect 307312 139534 307340 139567
rect 307300 139528 307352 139534
rect 307300 139470 307352 139476
rect 307298 138272 307354 138281
rect 307298 138207 307354 138216
rect 307312 138174 307340 138207
rect 307300 138168 307352 138174
rect 307300 138110 307352 138116
rect 307220 137142 307340 137170
rect 307206 137048 307262 137057
rect 307206 136983 307262 136992
rect 307036 133334 307156 133362
rect 306564 132660 306616 132666
rect 306564 132602 306616 132608
rect 306562 132288 306618 132297
rect 306562 132223 306618 132232
rect 306576 131170 306604 132223
rect 306930 131880 306986 131889
rect 306930 131815 306986 131824
rect 306944 131238 306972 131815
rect 306932 131232 306984 131238
rect 306932 131174 306984 131180
rect 306564 131164 306616 131170
rect 306564 131106 306616 131112
rect 306562 126848 306618 126857
rect 306562 126783 306618 126792
rect 305736 126268 305788 126274
rect 305736 126210 305788 126216
rect 306576 125730 306604 126783
rect 306564 125724 306616 125730
rect 306564 125666 306616 125672
rect 306562 125488 306618 125497
rect 306562 125423 306618 125432
rect 306576 124370 306604 125423
rect 306564 124364 306616 124370
rect 306564 124306 306616 124312
rect 306562 118688 306618 118697
rect 306562 118623 306618 118632
rect 306576 117570 306604 118623
rect 306564 117564 306616 117570
rect 306564 117506 306616 117512
rect 306930 116648 306986 116657
rect 307036 116618 307064 133334
rect 307114 133240 307170 133249
rect 307114 133175 307170 133184
rect 307128 132598 307156 133175
rect 307116 132592 307168 132598
rect 307116 132534 307168 132540
rect 307114 121272 307170 121281
rect 307114 121207 307170 121216
rect 307128 120154 307156 121207
rect 307116 120148 307168 120154
rect 307116 120090 307168 120096
rect 307114 120048 307170 120057
rect 307114 119983 307170 119992
rect 307128 118726 307156 119983
rect 307116 118720 307168 118726
rect 307116 118662 307168 118668
rect 307114 117464 307170 117473
rect 307114 117399 307170 117408
rect 307128 117366 307156 117399
rect 307116 117360 307168 117366
rect 307116 117302 307168 117308
rect 306930 116583 306986 116592
rect 307024 116612 307076 116618
rect 306944 116074 306972 116583
rect 307024 116554 307076 116560
rect 307022 116240 307078 116249
rect 307022 116175 307078 116184
rect 306932 116068 306984 116074
rect 306932 116010 306984 116016
rect 305826 108080 305882 108089
rect 305826 108015 305882 108024
rect 305644 107636 305696 107642
rect 305644 107578 305696 107584
rect 304632 106344 304684 106350
rect 304632 106286 304684 106292
rect 304540 105596 304592 105602
rect 304540 105538 304592 105544
rect 304644 69698 304672 106286
rect 305642 105360 305698 105369
rect 305642 105295 305698 105304
rect 304632 69692 304684 69698
rect 304632 69634 304684 69640
rect 304448 54596 304500 54602
rect 304448 54538 304500 54544
rect 304356 25560 304408 25566
rect 304356 25502 304408 25508
rect 305656 6254 305684 105295
rect 305734 101144 305790 101153
rect 305734 101079 305790 101088
rect 305748 42090 305776 101079
rect 305840 65618 305868 108015
rect 306746 106856 306802 106865
rect 306746 106791 306802 106800
rect 305918 106448 305974 106457
rect 305918 106383 305974 106392
rect 305932 73846 305960 106383
rect 306760 106350 306788 106791
rect 306748 106344 306800 106350
rect 306748 106286 306800 106292
rect 306746 100056 306802 100065
rect 306746 99991 306802 100000
rect 306760 99550 306788 99991
rect 306748 99544 306800 99550
rect 306748 99486 306800 99492
rect 306930 97472 306986 97481
rect 306930 97407 306986 97416
rect 306944 96762 306972 97407
rect 306932 96756 306984 96762
rect 306932 96698 306984 96704
rect 306930 96248 306986 96257
rect 306930 96183 306986 96192
rect 306944 95266 306972 96183
rect 306932 95260 306984 95266
rect 306932 95202 306984 95208
rect 305920 73840 305972 73846
rect 305920 73782 305972 73788
rect 305828 65612 305880 65618
rect 305828 65554 305880 65560
rect 305736 42084 305788 42090
rect 305736 42026 305788 42032
rect 306380 14612 306432 14618
rect 306380 14554 306432 14560
rect 305644 6248 305696 6254
rect 305644 6190 305696 6196
rect 304354 3496 304410 3505
rect 304354 3431 304410 3440
rect 305550 3496 305606 3505
rect 305550 3431 305606 3440
rect 304264 2168 304316 2174
rect 304264 2110 304316 2116
rect 304368 480 304396 3431
rect 305564 480 305592 3431
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306392 354 306420 14554
rect 307036 8974 307064 116175
rect 307114 115696 307170 115705
rect 307114 115631 307170 115640
rect 307128 114578 307156 115631
rect 307116 114572 307168 114578
rect 307116 114514 307168 114520
rect 307114 98696 307170 98705
rect 307114 98631 307170 98640
rect 307128 29646 307156 98631
rect 307220 87650 307248 136983
rect 307312 130422 307340 137142
rect 307404 134570 307432 140791
rect 307666 140448 307722 140457
rect 307666 140383 307722 140392
rect 307680 139466 307708 140383
rect 307668 139460 307720 139466
rect 307668 139402 307720 139408
rect 307574 139088 307630 139097
rect 307574 139023 307630 139032
rect 307588 138038 307616 139023
rect 307666 138680 307722 138689
rect 307666 138615 307722 138624
rect 307680 138106 307708 138615
rect 307668 138100 307720 138106
rect 307668 138042 307720 138048
rect 307576 138032 307628 138038
rect 307576 137974 307628 137980
rect 307574 137864 307630 137873
rect 307574 137799 307630 137808
rect 307588 136746 307616 137799
rect 307666 137456 307722 137465
rect 307666 137391 307722 137400
rect 307576 136740 307628 136746
rect 307576 136682 307628 136688
rect 307680 136678 307708 137391
rect 307668 136672 307720 136678
rect 307482 136640 307538 136649
rect 307668 136614 307720 136620
rect 307482 136575 307538 136584
rect 307496 135386 307524 136575
rect 307574 136232 307630 136241
rect 307574 136167 307630 136176
rect 307484 135380 307536 135386
rect 307484 135322 307536 135328
rect 307588 135318 307616 136167
rect 307668 135448 307720 135454
rect 307668 135390 307720 135396
rect 307576 135312 307628 135318
rect 307680 135289 307708 135390
rect 307576 135254 307628 135260
rect 307666 135280 307722 135289
rect 307666 135215 307722 135224
rect 307392 134564 307444 134570
rect 307392 134506 307444 134512
rect 307666 134464 307722 134473
rect 307666 134399 307722 134408
rect 307680 133958 307708 134399
rect 307668 133952 307720 133958
rect 307668 133894 307720 133900
rect 307666 132696 307722 132705
rect 307666 132631 307722 132640
rect 307680 132530 307708 132631
rect 307668 132524 307720 132530
rect 307668 132466 307720 132472
rect 307482 131064 307538 131073
rect 307482 130999 307538 131008
rect 307300 130416 307352 130422
rect 307300 130358 307352 130364
rect 307496 129878 307524 130999
rect 307666 129976 307722 129985
rect 307666 129911 307722 129920
rect 307484 129872 307536 129878
rect 307298 129840 307354 129849
rect 307484 129814 307536 129820
rect 307680 129810 307708 129911
rect 307298 129775 307354 129784
rect 307668 129804 307720 129810
rect 307312 91798 307340 129775
rect 307668 129746 307720 129752
rect 307574 129296 307630 129305
rect 307574 129231 307630 129240
rect 307484 128512 307536 128518
rect 307482 128480 307484 128489
rect 307536 128480 307538 128489
rect 307588 128450 307616 129231
rect 307666 128888 307722 128897
rect 307666 128823 307722 128832
rect 307482 128415 307538 128424
rect 307576 128444 307628 128450
rect 307576 128386 307628 128392
rect 307680 128382 307708 128823
rect 307668 128376 307720 128382
rect 307668 128318 307720 128324
rect 307482 128072 307538 128081
rect 307482 128007 307538 128016
rect 307496 127022 307524 128007
rect 307574 127664 307630 127673
rect 307574 127599 307630 127608
rect 307588 127158 307616 127599
rect 307666 127256 307722 127265
rect 307666 127191 307722 127200
rect 307576 127152 307628 127158
rect 307576 127094 307628 127100
rect 307680 127090 307708 127191
rect 307668 127084 307720 127090
rect 307668 127026 307720 127032
rect 307484 127016 307536 127022
rect 307484 126958 307536 126964
rect 307666 125896 307722 125905
rect 307666 125831 307722 125840
rect 307680 125662 307708 125831
rect 307668 125656 307720 125662
rect 307668 125598 307720 125604
rect 307574 125080 307630 125089
rect 307574 125015 307630 125024
rect 307484 124296 307536 124302
rect 307482 124264 307484 124273
rect 307536 124264 307538 124273
rect 307588 124234 307616 125015
rect 307666 124672 307722 124681
rect 307666 124607 307722 124616
rect 307680 124438 307708 124607
rect 307668 124432 307720 124438
rect 307668 124374 307720 124380
rect 307482 124199 307538 124208
rect 307576 124228 307628 124234
rect 307576 124170 307628 124176
rect 307482 123856 307538 123865
rect 307482 123791 307538 123800
rect 307496 122942 307524 123791
rect 307574 123448 307630 123457
rect 307574 123383 307630 123392
rect 307484 122936 307536 122942
rect 307484 122878 307536 122884
rect 307588 122874 307616 123383
rect 307666 123040 307722 123049
rect 307666 122975 307668 122984
rect 307720 122975 307722 122984
rect 307668 122946 307720 122952
rect 307576 122868 307628 122874
rect 307576 122810 307628 122816
rect 307574 122496 307630 122505
rect 307574 122431 307630 122440
rect 307482 121680 307538 121689
rect 307482 121615 307484 121624
rect 307536 121615 307538 121624
rect 307484 121586 307536 121592
rect 307588 121582 307616 122431
rect 307666 122088 307722 122097
rect 307666 122023 307722 122032
rect 307576 121576 307628 121582
rect 307576 121518 307628 121524
rect 307680 121514 307708 122023
rect 307668 121508 307720 121514
rect 307668 121450 307720 121456
rect 307574 120864 307630 120873
rect 307574 120799 307630 120808
rect 307588 120222 307616 120799
rect 307666 120456 307722 120465
rect 307666 120391 307722 120400
rect 307680 120290 307708 120391
rect 307668 120284 307720 120290
rect 307668 120226 307720 120232
rect 307576 120216 307628 120222
rect 307576 120158 307628 120164
rect 307574 119640 307630 119649
rect 307574 119575 307630 119584
rect 307588 118794 307616 119575
rect 307666 119096 307722 119105
rect 307666 119031 307722 119040
rect 307680 118862 307708 119031
rect 307668 118856 307720 118862
rect 307668 118798 307720 118804
rect 307576 118788 307628 118794
rect 307576 118730 307628 118736
rect 307574 118280 307630 118289
rect 307574 118215 307630 118224
rect 307588 117434 307616 118215
rect 307666 117872 307722 117881
rect 307666 117807 307722 117816
rect 307680 117502 307708 117807
rect 307668 117496 307720 117502
rect 307668 117438 307720 117444
rect 307576 117428 307628 117434
rect 307576 117370 307628 117376
rect 307666 117056 307722 117065
rect 307666 116991 307722 117000
rect 307680 116006 307708 116991
rect 307668 116000 307720 116006
rect 307668 115942 307720 115948
rect 307574 115288 307630 115297
rect 307574 115223 307630 115232
rect 307588 114646 307616 115223
rect 307666 114880 307722 114889
rect 307666 114815 307722 114824
rect 307680 114714 307708 114815
rect 307668 114708 307720 114714
rect 307668 114650 307720 114656
rect 307576 114640 307628 114646
rect 307576 114582 307628 114588
rect 307482 114472 307538 114481
rect 307482 114407 307538 114416
rect 307496 113218 307524 114407
rect 307574 113656 307630 113665
rect 307574 113591 307630 113600
rect 307588 113354 307616 113591
rect 307576 113348 307628 113354
rect 307576 113290 307628 113296
rect 307668 113280 307720 113286
rect 307666 113248 307668 113257
rect 307720 113248 307722 113257
rect 307484 113212 307536 113218
rect 307666 113183 307722 113192
rect 307484 113154 307536 113160
rect 307666 112704 307722 112713
rect 307666 112639 307722 112648
rect 307574 112296 307630 112305
rect 307574 112231 307630 112240
rect 307588 111926 307616 112231
rect 307680 111994 307708 112639
rect 307668 111988 307720 111994
rect 307668 111930 307720 111936
rect 307576 111920 307628 111926
rect 307576 111862 307628 111868
rect 307666 111888 307722 111897
rect 307666 111823 307668 111832
rect 307720 111823 307722 111832
rect 307668 111794 307720 111800
rect 307574 111480 307630 111489
rect 307574 111415 307630 111424
rect 307482 111072 307538 111081
rect 307482 111007 307538 111016
rect 307496 110634 307524 111007
rect 307484 110628 307536 110634
rect 307484 110570 307536 110576
rect 307588 110498 307616 111415
rect 307666 110664 307722 110673
rect 307666 110599 307722 110608
rect 307680 110566 307708 110599
rect 307668 110560 307720 110566
rect 307668 110502 307720 110508
rect 307576 110492 307628 110498
rect 307576 110434 307628 110440
rect 307482 110256 307538 110265
rect 307482 110191 307538 110200
rect 307496 109206 307524 110191
rect 307574 109848 307630 109857
rect 307574 109783 307630 109792
rect 307484 109200 307536 109206
rect 307484 109142 307536 109148
rect 307588 109138 307616 109783
rect 307666 109304 307722 109313
rect 307666 109239 307722 109248
rect 307576 109132 307628 109138
rect 307576 109074 307628 109080
rect 307680 109070 307708 109239
rect 307668 109064 307720 109070
rect 307668 109006 307720 109012
rect 307666 108896 307722 108905
rect 307666 108831 307722 108840
rect 307574 108488 307630 108497
rect 307574 108423 307630 108432
rect 307484 107772 307536 107778
rect 307484 107714 307536 107720
rect 307496 107681 307524 107714
rect 307588 107710 307616 108423
rect 307680 107914 307708 108831
rect 307668 107908 307720 107914
rect 307668 107850 307720 107856
rect 307576 107704 307628 107710
rect 307482 107672 307538 107681
rect 307576 107646 307628 107652
rect 307482 107607 307538 107616
rect 307666 107264 307722 107273
rect 307666 107199 307722 107208
rect 307680 106418 307708 107199
rect 307668 106412 307720 106418
rect 307668 106354 307720 106360
rect 307574 105904 307630 105913
rect 307574 105839 307630 105848
rect 307588 104922 307616 105839
rect 307666 105088 307722 105097
rect 307666 105023 307668 105032
rect 307720 105023 307722 105032
rect 307668 104994 307720 105000
rect 307576 104916 307628 104922
rect 307576 104858 307628 104864
rect 307482 104680 307538 104689
rect 307482 104615 307538 104624
rect 307496 103698 307524 104615
rect 307574 104272 307630 104281
rect 307574 104207 307630 104216
rect 307484 103692 307536 103698
rect 307484 103634 307536 103640
rect 307588 103630 307616 104207
rect 307666 103864 307722 103873
rect 307666 103799 307722 103808
rect 307576 103624 307628 103630
rect 307576 103566 307628 103572
rect 307680 103562 307708 103799
rect 307668 103556 307720 103562
rect 307668 103498 307720 103504
rect 307482 103456 307538 103465
rect 307482 103391 307538 103400
rect 307496 102202 307524 103391
rect 307574 103048 307630 103057
rect 307574 102983 307630 102992
rect 307588 102338 307616 102983
rect 307666 102504 307722 102513
rect 307666 102439 307722 102448
rect 307576 102332 307628 102338
rect 307576 102274 307628 102280
rect 307680 102270 307708 102439
rect 307668 102264 307720 102270
rect 307668 102206 307720 102212
rect 307484 102196 307536 102202
rect 307484 102138 307536 102144
rect 307574 102096 307630 102105
rect 307574 102031 307630 102040
rect 307482 101008 307538 101017
rect 307588 100978 307616 102031
rect 307482 100943 307538 100952
rect 307576 100972 307628 100978
rect 307496 100842 307524 100943
rect 307576 100914 307628 100920
rect 307668 100904 307720 100910
rect 307666 100872 307668 100881
rect 307720 100872 307722 100881
rect 307484 100836 307536 100842
rect 307666 100807 307722 100816
rect 307484 100778 307536 100784
rect 307574 100464 307630 100473
rect 307574 100399 307630 100408
rect 307588 99414 307616 100399
rect 307666 99648 307722 99657
rect 307666 99583 307722 99592
rect 307680 99482 307708 99583
rect 307668 99476 307720 99482
rect 307668 99418 307720 99424
rect 307576 99408 307628 99414
rect 307576 99350 307628 99356
rect 307574 99104 307630 99113
rect 307574 99039 307630 99048
rect 307588 98122 307616 99039
rect 307666 98288 307722 98297
rect 307666 98223 307722 98232
rect 307576 98116 307628 98122
rect 307576 98058 307628 98064
rect 307680 98054 307708 98223
rect 307668 98048 307720 98054
rect 307668 97990 307720 97996
rect 307666 97880 307722 97889
rect 307666 97815 307722 97824
rect 307680 96830 307708 97815
rect 307668 96824 307720 96830
rect 307668 96766 307720 96772
rect 307668 96688 307720 96694
rect 307666 96656 307668 96665
rect 307720 96656 307722 96665
rect 307666 96591 307722 96600
rect 307300 91792 307352 91798
rect 307300 91734 307352 91740
rect 307208 87644 307260 87650
rect 307208 87586 307260 87592
rect 307760 86284 307812 86290
rect 307760 86226 307812 86232
rect 307116 29640 307168 29646
rect 307116 29582 307168 29588
rect 307024 8968 307076 8974
rect 307024 8910 307076 8916
rect 307772 3482 307800 86226
rect 307850 30968 307906 30977
rect 307850 30903 307906 30912
rect 307864 3602 307892 30903
rect 308416 3670 308444 322186
rect 308496 265056 308548 265062
rect 308496 264998 308548 265004
rect 308508 95062 308536 264998
rect 308586 134872 308642 134881
rect 308586 134807 308642 134816
rect 308496 95056 308548 95062
rect 308496 94998 308548 95004
rect 308600 35222 308628 134807
rect 308588 35216 308640 35222
rect 308588 35158 308640 35164
rect 309140 21548 309192 21554
rect 309140 21490 309192 21496
rect 309152 16574 309180 21490
rect 309152 16546 309640 16574
rect 308404 3664 308456 3670
rect 308404 3606 308456 3612
rect 307852 3596 307904 3602
rect 307852 3538 307904 3544
rect 309048 3596 309100 3602
rect 309048 3538 309100 3544
rect 307772 3454 307984 3482
rect 307956 480 307984 3454
rect 309060 480 309088 3538
rect 309612 490 309640 16546
rect 309796 6914 309824 385018
rect 309876 334620 309928 334626
rect 309876 334562 309928 334568
rect 309704 6886 309824 6914
rect 309704 4146 309732 6886
rect 309692 4140 309744 4146
rect 309692 4082 309744 4088
rect 309888 3602 309916 334562
rect 311164 284368 311216 284374
rect 311164 284310 311216 284316
rect 311176 183054 311204 284310
rect 312544 278792 312596 278798
rect 312544 278734 312596 278740
rect 311256 220176 311308 220182
rect 311256 220118 311308 220124
rect 311164 183048 311216 183054
rect 311164 182990 311216 182996
rect 311268 178770 311296 220118
rect 311256 178764 311308 178770
rect 311256 178706 311308 178712
rect 312556 176118 312584 278734
rect 313936 177449 313964 386378
rect 324964 367124 325016 367130
rect 324964 367066 325016 367072
rect 316776 364404 316828 364410
rect 316776 364346 316828 364352
rect 316684 343664 316736 343670
rect 316684 343606 316736 343612
rect 315304 277500 315356 277506
rect 315304 277442 315356 277448
rect 314016 253972 314068 253978
rect 314016 253914 314068 253920
rect 314028 177478 314056 253914
rect 315316 178838 315344 277442
rect 316696 253201 316724 343606
rect 316788 339454 316816 364346
rect 316776 339448 316828 339454
rect 316776 339390 316828 339396
rect 319444 302320 319496 302326
rect 319444 302262 319496 302268
rect 318064 298308 318116 298314
rect 318064 298250 318116 298256
rect 316682 253192 316738 253201
rect 316682 253127 316738 253136
rect 316684 213240 316736 213246
rect 316684 213182 316736 213188
rect 315304 178832 315356 178838
rect 315304 178774 315356 178780
rect 316040 178084 316092 178090
rect 316040 178026 316092 178032
rect 314016 177472 314068 177478
rect 313922 177440 313978 177449
rect 314016 177414 314068 177420
rect 313922 177375 313978 177384
rect 312544 176112 312596 176118
rect 312544 176054 312596 176060
rect 316052 175930 316080 178026
rect 316696 176050 316724 213182
rect 316684 176044 316736 176050
rect 316684 175986 316736 175992
rect 318076 175982 318104 298250
rect 319456 176186 319484 302262
rect 320824 298172 320876 298178
rect 320824 298114 320876 298120
rect 319536 295384 319588 295390
rect 319536 295326 319588 295332
rect 319548 177614 319576 295326
rect 319628 188488 319680 188494
rect 319628 188430 319680 188436
rect 319536 177608 319588 177614
rect 319536 177550 319588 177556
rect 319640 177546 319668 188430
rect 319628 177540 319680 177546
rect 319628 177482 319680 177488
rect 319444 176180 319496 176186
rect 319444 176122 319496 176128
rect 316020 175902 316080 175930
rect 318064 175976 318116 175982
rect 320836 175953 320864 298114
rect 322204 277432 322256 277438
rect 322204 277374 322256 277380
rect 321560 243568 321612 243574
rect 321560 243510 321612 243516
rect 320916 233980 320968 233986
rect 320916 233922 320968 233928
rect 320928 190454 320956 233922
rect 320928 190426 321324 190454
rect 318064 175918 318116 175924
rect 320822 175944 320878 175953
rect 320822 175879 320878 175888
rect 321296 169697 321324 190426
rect 321468 176112 321520 176118
rect 321468 176054 321520 176060
rect 321480 175273 321508 176054
rect 321466 175264 321522 175273
rect 321466 175199 321522 175208
rect 321282 169688 321338 169697
rect 321282 169623 321338 169632
rect 321572 119921 321600 243510
rect 321744 192500 321796 192506
rect 321744 192442 321796 192448
rect 321652 182844 321704 182850
rect 321652 182786 321704 182792
rect 321664 127537 321692 182786
rect 321756 159905 321784 192442
rect 321742 159896 321798 159905
rect 321742 159831 321798 159840
rect 322216 142390 322244 277374
rect 324976 236706 325004 367066
rect 341536 333946 341564 700266
rect 397472 699718 397500 703520
rect 413664 702982 413692 703520
rect 413652 702976 413704 702982
rect 413652 702918 413704 702924
rect 429856 702846 429884 703520
rect 462332 702914 462360 703520
rect 462320 702908 462372 702914
rect 462320 702850 462372 702856
rect 429844 702840 429896 702846
rect 429844 702782 429896 702788
rect 478524 702778 478552 703520
rect 478512 702772 478564 702778
rect 478512 702714 478564 702720
rect 494808 702710 494836 703520
rect 494796 702704 494848 702710
rect 494796 702646 494848 702652
rect 527192 702574 527220 703520
rect 527180 702568 527232 702574
rect 527180 702510 527232 702516
rect 543476 702506 543504 703520
rect 559668 702642 559696 703520
rect 559656 702636 559708 702642
rect 559656 702578 559708 702584
rect 543464 702500 543516 702506
rect 543464 702442 543516 702448
rect 395344 699712 395396 699718
rect 395344 699654 395396 699660
rect 397460 699712 397512 699718
rect 397460 699654 397512 699660
rect 353300 389224 353352 389230
rect 353300 389166 353352 389172
rect 349160 373312 349212 373318
rect 349160 373254 349212 373260
rect 346400 348424 346452 348430
rect 346400 348366 346452 348372
rect 343640 336116 343692 336122
rect 343640 336058 343692 336064
rect 341524 333940 341576 333946
rect 341524 333882 341576 333888
rect 333244 299600 333296 299606
rect 333244 299542 333296 299548
rect 328736 286340 328788 286346
rect 328736 286282 328788 286288
rect 325700 282940 325752 282946
rect 325700 282882 325752 282888
rect 324964 236700 325016 236706
rect 324964 236642 325016 236648
rect 324594 217288 324650 217297
rect 324594 217223 324650 217232
rect 322940 215960 322992 215966
rect 322940 215902 322992 215908
rect 322204 142384 322256 142390
rect 322204 142326 322256 142332
rect 321650 127528 321706 127537
rect 321650 127463 321706 127472
rect 322952 120873 322980 215902
rect 323124 186992 323176 186998
rect 323124 186934 323176 186940
rect 323030 181384 323086 181393
rect 323030 181319 323086 181328
rect 323044 121689 323072 181319
rect 323136 150929 323164 186934
rect 324320 185632 324372 185638
rect 324320 185574 324372 185580
rect 323216 184272 323268 184278
rect 323216 184214 323268 184220
rect 323228 170105 323256 184214
rect 324332 174049 324360 185574
rect 324412 177336 324464 177342
rect 324412 177278 324464 177284
rect 324318 174040 324374 174049
rect 324318 173975 324374 173984
rect 324320 173868 324372 173874
rect 324320 173810 324372 173816
rect 324332 173233 324360 173810
rect 324318 173224 324374 173233
rect 324318 173159 324374 173168
rect 324424 172417 324452 177278
rect 324410 172408 324466 172417
rect 324410 172343 324466 172352
rect 324320 171080 324372 171086
rect 324320 171022 324372 171028
rect 324332 170921 324360 171022
rect 324318 170912 324374 170921
rect 324318 170847 324374 170856
rect 323214 170096 323270 170105
rect 323214 170031 323270 170040
rect 324320 169720 324372 169726
rect 324320 169662 324372 169668
rect 324332 168609 324360 169662
rect 324318 168600 324374 168609
rect 324318 168535 324374 168544
rect 324320 168360 324372 168366
rect 324320 168302 324372 168308
rect 324332 167793 324360 168302
rect 324412 168292 324464 168298
rect 324412 168234 324464 168240
rect 324318 167784 324374 167793
rect 324318 167719 324374 167728
rect 324424 167113 324452 168234
rect 324410 167104 324466 167113
rect 324410 167039 324466 167048
rect 324320 167000 324372 167006
rect 324320 166942 324372 166948
rect 324332 166297 324360 166942
rect 324318 166288 324374 166297
rect 324318 166223 324374 166232
rect 324412 165572 324464 165578
rect 324412 165514 324464 165520
rect 324320 165504 324372 165510
rect 324318 165472 324320 165481
rect 324372 165472 324374 165481
rect 324318 165407 324374 165416
rect 324424 164801 324452 165514
rect 324410 164792 324466 164801
rect 324410 164727 324466 164736
rect 324412 164212 324464 164218
rect 324412 164154 324464 164160
rect 324320 164144 324372 164150
rect 324320 164086 324372 164092
rect 324332 163985 324360 164086
rect 324318 163976 324374 163985
rect 324318 163911 324374 163920
rect 324424 163169 324452 164154
rect 324410 163160 324466 163169
rect 324410 163095 324466 163104
rect 324412 162852 324464 162858
rect 324412 162794 324464 162800
rect 324320 162784 324372 162790
rect 324320 162726 324372 162732
rect 324332 162489 324360 162726
rect 324318 162480 324374 162489
rect 324318 162415 324374 162424
rect 324424 161673 324452 162794
rect 324410 161664 324466 161673
rect 324410 161599 324466 161608
rect 324320 161424 324372 161430
rect 324320 161366 324372 161372
rect 324332 160857 324360 161366
rect 324412 161356 324464 161362
rect 324412 161298 324464 161304
rect 324318 160848 324374 160857
rect 324318 160783 324374 160792
rect 324424 160177 324452 161298
rect 324410 160168 324466 160177
rect 324410 160103 324466 160112
rect 324412 158704 324464 158710
rect 324412 158646 324464 158652
rect 324320 158636 324372 158642
rect 324320 158578 324372 158584
rect 324332 158545 324360 158578
rect 324318 158536 324374 158545
rect 324318 158471 324374 158480
rect 324424 157865 324452 158646
rect 324410 157856 324466 157865
rect 324410 157791 324466 157800
rect 324320 157276 324372 157282
rect 324320 157218 324372 157224
rect 324332 157049 324360 157218
rect 324318 157040 324374 157049
rect 324318 156975 324374 156984
rect 324320 156868 324372 156874
rect 324320 156810 324372 156816
rect 324332 156369 324360 156810
rect 324318 156360 324374 156369
rect 324318 156295 324374 156304
rect 324412 155916 324464 155922
rect 324412 155858 324464 155864
rect 324320 155848 324372 155854
rect 324320 155790 324372 155796
rect 324332 155553 324360 155790
rect 324318 155544 324374 155553
rect 324318 155479 324374 155488
rect 324424 154737 324452 155858
rect 324410 154728 324466 154737
rect 324410 154663 324466 154672
rect 324320 154556 324372 154562
rect 324320 154498 324372 154504
rect 324332 154057 324360 154498
rect 324318 154048 324374 154057
rect 324318 153983 324374 153992
rect 324320 153468 324372 153474
rect 324320 153410 324372 153416
rect 324332 153241 324360 153410
rect 324318 153232 324374 153241
rect 324318 153167 324374 153176
rect 324412 153196 324464 153202
rect 324412 153138 324464 153144
rect 324424 152425 324452 153138
rect 324410 152416 324466 152425
rect 324410 152351 324466 152360
rect 324320 151768 324372 151774
rect 324318 151736 324320 151745
rect 324372 151736 324374 151745
rect 324318 151671 324374 151680
rect 323122 150920 323178 150929
rect 323122 150855 323178 150864
rect 324320 150408 324372 150414
rect 324320 150350 324372 150356
rect 324332 150113 324360 150350
rect 324412 150340 324464 150346
rect 324412 150282 324464 150288
rect 324318 150104 324374 150113
rect 324318 150039 324374 150048
rect 324424 149433 324452 150282
rect 324410 149424 324466 149433
rect 324410 149359 324466 149368
rect 324320 148980 324372 148986
rect 324320 148922 324372 148928
rect 324332 148617 324360 148922
rect 324318 148608 324374 148617
rect 324318 148543 324374 148552
rect 324320 147620 324372 147626
rect 324320 147562 324372 147568
rect 324332 147121 324360 147562
rect 324318 147112 324374 147121
rect 324318 147047 324374 147056
rect 324318 146296 324374 146305
rect 324318 146231 324320 146240
rect 324372 146231 324374 146240
rect 324320 146202 324372 146208
rect 324320 145716 324372 145722
rect 324320 145658 324372 145664
rect 324332 145489 324360 145658
rect 324318 145480 324374 145489
rect 324318 145415 324374 145424
rect 324412 144900 324464 144906
rect 324412 144842 324464 144848
rect 324320 144832 324372 144838
rect 324318 144800 324320 144809
rect 324372 144800 324374 144809
rect 324318 144735 324374 144744
rect 324424 143993 324452 144842
rect 324410 143984 324466 143993
rect 324410 143919 324466 143928
rect 324412 143540 324464 143546
rect 324412 143482 324464 143488
rect 324320 143472 324372 143478
rect 324320 143414 324372 143420
rect 324332 143177 324360 143414
rect 324318 143168 324374 143177
rect 324318 143103 324374 143112
rect 324424 142497 324452 143482
rect 324410 142488 324466 142497
rect 324410 142423 324466 142432
rect 324412 142384 324464 142390
rect 324412 142326 324464 142332
rect 324320 142044 324372 142050
rect 324320 141986 324372 141992
rect 324332 141681 324360 141986
rect 324318 141672 324374 141681
rect 324318 141607 324374 141616
rect 324320 140752 324372 140758
rect 324320 140694 324372 140700
rect 324332 140185 324360 140694
rect 324318 140176 324374 140185
rect 324318 140111 324374 140120
rect 324320 139392 324372 139398
rect 324318 139360 324320 139369
rect 324372 139360 324374 139369
rect 324318 139295 324374 139304
rect 324320 137896 324372 137902
rect 324318 137864 324320 137873
rect 324372 137864 324374 137873
rect 324318 137799 324374 137808
rect 324320 136400 324372 136406
rect 324318 136368 324320 136377
rect 324372 136368 324374 136377
rect 324318 136303 324374 136312
rect 324320 135244 324372 135250
rect 324320 135186 324372 135192
rect 324332 134745 324360 135186
rect 324318 134736 324374 134745
rect 324318 134671 324374 134680
rect 324320 133884 324372 133890
rect 324320 133826 324372 133832
rect 324332 133249 324360 133826
rect 324318 133240 324374 133249
rect 324318 133175 324374 133184
rect 324424 132494 324452 142326
rect 324504 142112 324556 142118
rect 324504 142054 324556 142060
rect 324516 140865 324544 142054
rect 324502 140856 324558 140865
rect 324502 140791 324558 140800
rect 324504 139324 324556 139330
rect 324504 139266 324556 139272
rect 324516 138553 324544 139266
rect 324502 138544 324558 138553
rect 324502 138479 324558 138488
rect 324504 137964 324556 137970
rect 324504 137906 324556 137912
rect 324516 137057 324544 137906
rect 324502 137048 324558 137057
rect 324502 136983 324558 136992
rect 324504 136604 324556 136610
rect 324504 136546 324556 136552
rect 324516 135561 324544 136546
rect 324502 135552 324558 135561
rect 324502 135487 324558 135496
rect 324424 132466 324544 132494
rect 324320 131096 324372 131102
rect 324320 131038 324372 131044
rect 324332 130937 324360 131038
rect 324412 131028 324464 131034
rect 324412 130970 324464 130976
rect 324318 130928 324374 130937
rect 324318 130863 324374 130872
rect 324424 130121 324452 130970
rect 324410 130112 324466 130121
rect 324410 130047 324466 130056
rect 324320 129736 324372 129742
rect 324320 129678 324372 129684
rect 324332 129441 324360 129678
rect 324412 129668 324464 129674
rect 324412 129610 324464 129616
rect 324318 129432 324374 129441
rect 324318 129367 324374 129376
rect 324424 128625 324452 129610
rect 324410 128616 324466 128625
rect 324410 128551 324466 128560
rect 324320 128308 324372 128314
rect 324320 128250 324372 128256
rect 324332 127809 324360 128250
rect 324318 127800 324374 127809
rect 324318 127735 324374 127744
rect 324516 126313 324544 132466
rect 324502 126304 324558 126313
rect 324502 126239 324558 126248
rect 324320 125588 324372 125594
rect 324320 125530 324372 125536
rect 324332 125497 324360 125530
rect 324318 125488 324374 125497
rect 324318 125423 324374 125432
rect 324320 124160 324372 124166
rect 324320 124102 324372 124108
rect 324332 124001 324360 124102
rect 324412 124092 324464 124098
rect 324412 124034 324464 124040
rect 324318 123992 324374 124001
rect 324318 123927 324374 123936
rect 324424 123185 324452 124034
rect 324410 123176 324466 123185
rect 324410 123111 324466 123120
rect 324320 122800 324372 122806
rect 324320 122742 324372 122748
rect 324332 122505 324360 122742
rect 324318 122496 324374 122505
rect 324318 122431 324374 122440
rect 323030 121680 323086 121689
rect 323030 121615 323086 121624
rect 324320 121440 324372 121446
rect 324320 121382 324372 121388
rect 322938 120864 322994 120873
rect 322938 120799 322994 120808
rect 324332 120193 324360 121382
rect 324318 120184 324374 120193
rect 324318 120119 324374 120128
rect 321558 119912 321614 119921
rect 321558 119847 321614 119856
rect 324412 118652 324464 118658
rect 324412 118594 324464 118600
rect 324320 118584 324372 118590
rect 324318 118552 324320 118561
rect 324372 118552 324374 118561
rect 324318 118487 324374 118496
rect 324424 117881 324452 118594
rect 324410 117872 324466 117881
rect 324410 117807 324466 117816
rect 324320 117292 324372 117298
rect 324320 117234 324372 117240
rect 324332 116385 324360 117234
rect 324318 116376 324374 116385
rect 324318 116311 324374 116320
rect 324412 115932 324464 115938
rect 324412 115874 324464 115880
rect 324320 115864 324372 115870
rect 324320 115806 324372 115812
rect 324332 115569 324360 115806
rect 324318 115560 324374 115569
rect 324318 115495 324374 115504
rect 324424 114753 324452 115874
rect 324410 114744 324466 114753
rect 324410 114679 324466 114688
rect 324412 114504 324464 114510
rect 324412 114446 324464 114452
rect 324320 114436 324372 114442
rect 324320 114378 324372 114384
rect 324332 114073 324360 114378
rect 324318 114064 324374 114073
rect 324318 113999 324374 114008
rect 324424 113257 324452 114446
rect 324410 113248 324466 113257
rect 324410 113183 324466 113192
rect 324320 113144 324372 113150
rect 324320 113086 324372 113092
rect 324332 112441 324360 113086
rect 324318 112432 324374 112441
rect 324318 112367 324374 112376
rect 324320 111784 324372 111790
rect 324320 111726 324372 111732
rect 324332 110945 324360 111726
rect 324318 110936 324374 110945
rect 324318 110871 324374 110880
rect 324412 110424 324464 110430
rect 324412 110366 324464 110372
rect 324320 110356 324372 110362
rect 324320 110298 324372 110304
rect 324332 110129 324360 110298
rect 324318 110120 324374 110129
rect 324318 110055 324374 110064
rect 324424 109449 324452 110366
rect 324410 109440 324466 109449
rect 324410 109375 324466 109384
rect 324320 108996 324372 109002
rect 324320 108938 324372 108944
rect 324332 107817 324360 108938
rect 324410 108624 324466 108633
rect 324410 108559 324466 108568
rect 324318 107808 324374 107817
rect 324318 107743 324374 107752
rect 324320 106276 324372 106282
rect 324320 106218 324372 106224
rect 324332 105505 324360 106218
rect 324318 105496 324374 105505
rect 324318 105431 324374 105440
rect 324318 104816 324374 104825
rect 324318 104751 324374 104760
rect 324332 103358 324360 104751
rect 324320 103352 324372 103358
rect 324320 103294 324372 103300
rect 324320 103216 324372 103222
rect 324318 103184 324320 103193
rect 324372 103184 324374 103193
rect 324318 103119 324374 103128
rect 324320 100700 324372 100706
rect 324320 100642 324372 100648
rect 321282 100464 321338 100473
rect 321282 100399 321338 100408
rect 321296 96626 321324 100399
rect 324332 100201 324360 100642
rect 324318 100192 324374 100201
rect 324318 100127 324374 100136
rect 321374 98832 321430 98841
rect 321374 98767 321430 98776
rect 321284 96620 321336 96626
rect 321284 96562 321336 96568
rect 321388 95169 321416 98767
rect 321558 97336 321614 97345
rect 321558 97271 321614 97280
rect 321466 96656 321522 96665
rect 321466 96591 321522 96600
rect 321480 96558 321508 96591
rect 321468 96552 321520 96558
rect 321468 96494 321520 96500
rect 321374 95160 321430 95169
rect 321374 95095 321430 95104
rect 321572 95062 321600 97271
rect 324424 95198 324452 108559
rect 324504 103488 324556 103494
rect 324504 103430 324556 103436
rect 324516 102513 324544 103430
rect 324502 102504 324558 102513
rect 324502 102439 324558 102448
rect 324608 98569 324636 217223
rect 325712 142186 325740 282882
rect 327172 238060 327224 238066
rect 327172 238002 327224 238008
rect 325792 218748 325844 218754
rect 325792 218690 325844 218696
rect 324964 142180 325016 142186
rect 324964 142122 325016 142128
rect 325700 142180 325752 142186
rect 325700 142122 325752 142128
rect 324976 132433 325004 142122
rect 324962 132424 325018 132433
rect 324962 132359 325018 132368
rect 325606 104000 325662 104009
rect 325804 103986 325832 218690
rect 327080 213308 327132 213314
rect 327080 213250 327132 213256
rect 325976 185836 326028 185842
rect 325976 185778 326028 185784
rect 325884 182912 325936 182918
rect 325884 182854 325936 182860
rect 325896 147801 325924 182854
rect 325988 156874 326016 185778
rect 326160 176180 326212 176186
rect 326160 176122 326212 176128
rect 326066 175944 326122 175953
rect 326066 175879 326122 175888
rect 326080 171193 326108 175879
rect 326172 173874 326200 176122
rect 326160 173868 326212 173874
rect 326160 173810 326212 173816
rect 326066 171184 326122 171193
rect 326066 171119 326122 171128
rect 325976 156868 326028 156874
rect 325976 156810 326028 156816
rect 325882 147792 325938 147801
rect 325882 147727 325938 147736
rect 325662 103958 325832 103986
rect 325606 103935 325662 103944
rect 324688 103352 324740 103358
rect 324688 103294 324740 103300
rect 324594 98560 324650 98569
rect 324594 98495 324650 98504
rect 324412 95192 324464 95198
rect 324412 95134 324464 95140
rect 324700 95130 324728 103294
rect 327092 103222 327120 213250
rect 327184 145722 327212 238002
rect 328644 200796 328696 200802
rect 328644 200738 328696 200744
rect 328552 196648 328604 196654
rect 328552 196590 328604 196596
rect 327356 185700 327408 185706
rect 327356 185642 327408 185648
rect 327264 180124 327316 180130
rect 327264 180066 327316 180072
rect 327172 145716 327224 145722
rect 327172 145658 327224 145664
rect 327276 136406 327304 180066
rect 327368 153474 327396 185642
rect 327356 153468 327408 153474
rect 327356 153410 327408 153416
rect 327264 136400 327316 136406
rect 327264 136342 327316 136348
rect 328564 128314 328592 196590
rect 328656 151774 328684 200738
rect 328644 151768 328696 151774
rect 328644 151710 328696 151716
rect 328748 140758 328776 286282
rect 331312 251252 331364 251258
rect 331312 251194 331364 251200
rect 329840 240168 329892 240174
rect 329840 240110 329892 240116
rect 328736 140752 328788 140758
rect 328736 140694 328788 140700
rect 329852 129674 329880 240110
rect 329932 199436 329984 199442
rect 329932 199378 329984 199384
rect 329944 129742 329972 199378
rect 330024 198076 330076 198082
rect 330024 198018 330076 198024
rect 330036 131034 330064 198018
rect 330116 177608 330168 177614
rect 330116 177550 330168 177556
rect 330128 162790 330156 177550
rect 331220 177540 331272 177546
rect 331220 177482 331272 177488
rect 331232 168298 331260 177482
rect 331220 168292 331272 168298
rect 331220 168234 331272 168240
rect 330116 162784 330168 162790
rect 330116 162726 330168 162732
rect 331324 150346 331352 251194
rect 331496 211812 331548 211818
rect 331496 211754 331548 211760
rect 331404 191276 331456 191282
rect 331404 191218 331456 191224
rect 331312 150340 331364 150346
rect 331312 150282 331364 150288
rect 331416 135250 331444 191218
rect 331404 135244 331456 135250
rect 331404 135186 331456 135192
rect 330024 131028 330076 131034
rect 330024 130970 330076 130976
rect 329932 129736 329984 129742
rect 329932 129678 329984 129684
rect 329840 129668 329892 129674
rect 329840 129610 329892 129616
rect 328552 128308 328604 128314
rect 328552 128250 328604 128256
rect 327080 103216 327132 103222
rect 327080 103158 327132 103164
rect 331508 100706 331536 211754
rect 332784 183048 332836 183054
rect 332784 182990 332836 182996
rect 332600 180192 332652 180198
rect 332600 180134 332652 180140
rect 332612 110362 332640 180134
rect 332692 177472 332744 177478
rect 332692 177414 332744 177420
rect 332704 125594 332732 177414
rect 332796 161362 332824 182990
rect 333256 177342 333284 299542
rect 335360 299532 335412 299538
rect 335360 299474 335412 299480
rect 334072 266484 334124 266490
rect 334072 266426 334124 266432
rect 333980 228472 334032 228478
rect 333980 228414 334032 228420
rect 333244 177336 333296 177342
rect 333244 177278 333296 177284
rect 332876 176044 332928 176050
rect 332876 175986 332928 175992
rect 332888 164150 332916 175986
rect 332876 164144 332928 164150
rect 332876 164086 332928 164092
rect 332784 161356 332836 161362
rect 332784 161298 332836 161304
rect 332692 125588 332744 125594
rect 332692 125530 332744 125536
rect 333992 114442 334020 228414
rect 334084 158642 334112 266426
rect 334256 188352 334308 188358
rect 334256 188294 334308 188300
rect 334164 182980 334216 182986
rect 334164 182922 334216 182928
rect 334072 158636 334124 158642
rect 334072 158578 334124 158584
rect 334176 137902 334204 182922
rect 334268 150414 334296 188294
rect 334256 150408 334308 150414
rect 334256 150350 334308 150356
rect 335372 147626 335400 299474
rect 342258 298344 342314 298353
rect 342258 298279 342314 298288
rect 338212 276072 338264 276078
rect 338212 276014 338264 276020
rect 335544 242956 335596 242962
rect 335544 242898 335596 242904
rect 335452 210452 335504 210458
rect 335452 210394 335504 210400
rect 335360 147620 335412 147626
rect 335360 147562 335412 147568
rect 334164 137896 334216 137902
rect 334164 137838 334216 137844
rect 335464 114510 335492 210394
rect 335556 162858 335584 242898
rect 336740 229764 336792 229770
rect 336740 229706 336792 229712
rect 335636 193860 335688 193866
rect 335636 193802 335688 193808
rect 335544 162852 335596 162858
rect 335544 162794 335596 162800
rect 335648 137970 335676 193802
rect 336752 144838 336780 229706
rect 336832 189780 336884 189786
rect 336832 189722 336884 189728
rect 336740 144832 336792 144838
rect 336740 144774 336792 144780
rect 335636 137964 335688 137970
rect 335636 137906 335688 137912
rect 335452 114504 335504 114510
rect 335452 114446 335504 114452
rect 333980 114436 334032 114442
rect 333980 114378 334032 114384
rect 336844 110430 336872 189722
rect 336924 181552 336976 181558
rect 336924 181494 336976 181500
rect 336936 164218 336964 181494
rect 338120 177336 338172 177342
rect 338120 177278 338172 177284
rect 337016 175976 337068 175982
rect 337016 175918 337068 175924
rect 336924 164212 336976 164218
rect 336924 164154 336976 164160
rect 337028 161430 337056 175918
rect 338132 171086 338160 177278
rect 338120 171080 338172 171086
rect 338120 171022 338172 171028
rect 337016 161424 337068 161430
rect 337016 161366 337068 161372
rect 338224 144906 338252 276014
rect 339500 267776 339552 267782
rect 339500 267718 339552 267724
rect 338396 262268 338448 262274
rect 338396 262210 338448 262216
rect 338304 209092 338356 209098
rect 338304 209034 338356 209040
rect 338212 144900 338264 144906
rect 338212 144842 338264 144848
rect 338316 117298 338344 209034
rect 338408 124098 338436 262210
rect 338396 124092 338448 124098
rect 338396 124034 338448 124040
rect 338304 117292 338356 117298
rect 338304 117234 338356 117240
rect 339512 113150 339540 267718
rect 339592 239488 339644 239494
rect 339592 239430 339644 239436
rect 339604 168366 339632 239430
rect 340880 221468 340932 221474
rect 340880 221410 340932 221416
rect 339684 185768 339736 185774
rect 339684 185710 339736 185716
rect 339592 168360 339644 168366
rect 339592 168302 339644 168308
rect 339696 118590 339724 185710
rect 339776 178832 339828 178838
rect 339776 178774 339828 178780
rect 339788 155854 339816 178774
rect 339776 155848 339828 155854
rect 339776 155790 339828 155796
rect 339684 118584 339736 118590
rect 339684 118526 339736 118532
rect 339500 113144 339552 113150
rect 339500 113086 339552 113092
rect 340892 111790 340920 221410
rect 340972 194064 341024 194070
rect 340972 194006 341024 194012
rect 340984 124166 341012 194006
rect 341156 188420 341208 188426
rect 341156 188362 341208 188368
rect 341064 184204 341116 184210
rect 341064 184146 341116 184152
rect 341076 139330 341104 184146
rect 341168 155922 341196 188362
rect 341156 155916 341208 155922
rect 341156 155858 341208 155864
rect 341064 139324 341116 139330
rect 341064 139266 341116 139272
rect 342272 136610 342300 298279
rect 342352 296812 342404 296818
rect 342352 296754 342404 296760
rect 342364 146266 342392 296754
rect 342444 244316 342496 244322
rect 342444 244258 342496 244264
rect 342456 242894 342484 244258
rect 342444 242888 342496 242894
rect 342444 242830 342496 242836
rect 342444 239420 342496 239426
rect 342444 239362 342496 239368
rect 342352 146260 342404 146266
rect 342352 146202 342404 146208
rect 342260 136604 342312 136610
rect 342260 136546 342312 136552
rect 340972 124160 341024 124166
rect 340972 124102 341024 124108
rect 342456 115870 342484 239362
rect 342536 178764 342588 178770
rect 342536 178706 342588 178712
rect 342444 115864 342496 115870
rect 342444 115806 342496 115812
rect 340880 111784 340932 111790
rect 340880 111726 340932 111732
rect 336832 110424 336884 110430
rect 336832 110366 336884 110372
rect 332600 110356 332652 110362
rect 332600 110298 332652 110304
rect 342548 109002 342576 178706
rect 342536 108996 342588 109002
rect 342536 108938 342588 108944
rect 331496 100700 331548 100706
rect 331496 100642 331548 100648
rect 324688 95124 324740 95130
rect 324688 95066 324740 95072
rect 321560 95056 321612 95062
rect 321560 94998 321612 95004
rect 324320 89004 324372 89010
rect 324320 88946 324372 88952
rect 314660 83496 314712 83502
rect 314660 83438 314712 83444
rect 313280 60104 313332 60110
rect 313280 60046 313332 60052
rect 313292 16574 313320 60046
rect 313292 16546 313872 16574
rect 309876 3596 309928 3602
rect 309876 3538 309928 3544
rect 312636 3528 312688 3534
rect 312636 3470 312688 3476
rect 311440 3460 311492 3466
rect 311440 3402 311492 3408
rect 306718 354 306830 480
rect 306392 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309612 462 309824 490
rect 311452 480 311480 3402
rect 312648 480 312676 3470
rect 313844 480 313872 16546
rect 309796 354 309824 462
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314672 354 314700 83438
rect 316040 78056 316092 78062
rect 316040 77998 316092 78004
rect 316052 3482 316080 77998
rect 321560 77988 321612 77994
rect 321560 77930 321612 77936
rect 316132 61464 316184 61470
rect 316132 61406 316184 61412
rect 316144 3670 316172 61406
rect 321572 16574 321600 77930
rect 321572 16546 322152 16574
rect 318524 4140 318576 4146
rect 318524 4082 318576 4088
rect 316132 3664 316184 3670
rect 316132 3606 316184 3612
rect 317328 3664 317380 3670
rect 317328 3606 317380 3612
rect 316052 3454 316264 3482
rect 316236 480 316264 3454
rect 317340 480 317368 3606
rect 318536 480 318564 4082
rect 320916 3732 320968 3738
rect 320916 3674 320968 3680
rect 319718 3496 319774 3505
rect 319718 3431 319774 3440
rect 319732 480 319760 3431
rect 320928 480 320956 3674
rect 322124 480 322152 16546
rect 322940 15972 322992 15978
rect 322940 15914 322992 15920
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 322952 354 322980 15914
rect 324332 3346 324360 88946
rect 324412 84856 324464 84862
rect 324412 84798 324464 84804
rect 324424 3534 324452 84798
rect 329840 82136 329892 82142
rect 329840 82078 329892 82084
rect 325700 80708 325752 80714
rect 325700 80650 325752 80656
rect 325712 16574 325740 80650
rect 329852 16574 329880 82078
rect 343652 16574 343680 336058
rect 343732 298240 343784 298246
rect 343732 298182 343784 298188
rect 343744 139398 343772 298182
rect 345020 287088 345072 287094
rect 345020 287030 345072 287036
rect 343916 202156 343968 202162
rect 343916 202098 343968 202104
rect 343822 182880 343878 182889
rect 343822 182815 343878 182824
rect 343836 143478 343864 182815
rect 343928 165510 343956 202098
rect 343916 165504 343968 165510
rect 343916 165446 343968 165452
rect 345032 143546 345060 287030
rect 345112 224256 345164 224262
rect 345112 224198 345164 224204
rect 345020 143540 345072 143546
rect 345020 143482 345072 143488
rect 343824 143472 343876 143478
rect 343824 143414 343876 143420
rect 343732 139392 343784 139398
rect 343732 139334 343784 139340
rect 345124 118658 345152 224198
rect 345204 195356 345256 195362
rect 345204 195298 345256 195304
rect 345216 133890 345244 195298
rect 345296 181484 345348 181490
rect 345296 181426 345348 181432
rect 345308 169726 345336 181426
rect 345296 169720 345348 169726
rect 345296 169662 345348 169668
rect 345204 133884 345256 133890
rect 345204 133826 345256 133832
rect 345112 118652 345164 118658
rect 345112 118594 345164 118600
rect 346412 16574 346440 348366
rect 347964 266416 348016 266422
rect 347964 266358 348016 266364
rect 346492 264988 346544 264994
rect 346492 264930 346544 264936
rect 346504 142050 346532 264930
rect 347872 258120 347924 258126
rect 347872 258062 347924 258068
rect 347780 236700 347832 236706
rect 347780 236642 347832 236648
rect 346584 178696 346636 178702
rect 346584 178638 346636 178644
rect 346674 178664 346730 178673
rect 346596 165578 346624 178638
rect 346674 178599 346730 178608
rect 346688 167006 346716 178599
rect 346676 167000 346728 167006
rect 346676 166942 346728 166948
rect 346584 165572 346636 165578
rect 346584 165514 346636 165520
rect 346492 142044 346544 142050
rect 346492 141986 346544 141992
rect 347792 16574 347820 236642
rect 347884 131102 347912 258062
rect 347976 148986 348004 266358
rect 347964 148980 348016 148986
rect 347964 148922 348016 148928
rect 347872 131096 347924 131102
rect 347872 131038 347924 131044
rect 325712 16546 326384 16574
rect 329852 16546 330432 16574
rect 343652 16546 344600 16574
rect 346412 16546 346992 16574
rect 347792 16546 348096 16574
rect 324412 3528 324464 3534
rect 324412 3470 324464 3476
rect 325608 3528 325660 3534
rect 325608 3470 325660 3476
rect 324332 3318 324452 3346
rect 324424 480 324452 3318
rect 325620 480 325648 3470
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 16546
rect 328000 11824 328052 11830
rect 328000 11766 328052 11772
rect 328012 480 328040 11766
rect 329196 3596 329248 3602
rect 329196 3538 329248 3544
rect 329208 480 329236 3538
rect 330404 480 330432 16546
rect 336278 4040 336334 4049
rect 336278 3975 336334 3984
rect 335082 3632 335138 3641
rect 335082 3567 335138 3576
rect 331586 3496 331642 3505
rect 331586 3431 331642 3440
rect 332690 3496 332746 3505
rect 332690 3431 332746 3440
rect 333886 3496 333942 3505
rect 333886 3431 333942 3440
rect 331600 480 331628 3431
rect 332704 480 332732 3431
rect 333900 480 333928 3431
rect 335096 480 335124 3567
rect 336292 480 336320 3975
rect 337474 3496 337530 3505
rect 337474 3431 337530 3440
rect 338670 3496 338726 3505
rect 338670 3431 338726 3440
rect 339866 3496 339922 3505
rect 339866 3431 339922 3440
rect 340970 3496 341026 3505
rect 343362 3496 343418 3505
rect 340970 3431 341026 3440
rect 342168 3460 342220 3466
rect 337488 480 337516 3431
rect 338684 480 338712 3431
rect 339880 480 339908 3431
rect 340984 480 341012 3431
rect 343362 3431 343418 3440
rect 342168 3402 342220 3408
rect 342180 480 342208 3402
rect 343376 480 343404 3431
rect 344572 480 344600 16546
rect 345754 3496 345810 3505
rect 345754 3431 345810 3440
rect 345768 480 345796 3431
rect 346964 480 346992 16546
rect 348068 480 348096 16546
rect 349172 3534 349200 373254
rect 349252 320884 349304 320890
rect 349252 320826 349304 320832
rect 349160 3528 349212 3534
rect 349160 3470 349212 3476
rect 349264 480 349292 320826
rect 349344 302252 349396 302258
rect 349344 302194 349396 302200
rect 349356 157282 349384 302194
rect 352010 295352 352066 295361
rect 352010 295287 352066 295296
rect 351920 292596 351972 292602
rect 351920 292538 351972 292544
rect 350632 291236 350684 291242
rect 350632 291178 350684 291184
rect 350540 177404 350592 177410
rect 350540 177346 350592 177352
rect 349344 157276 349396 157282
rect 349344 157218 349396 157224
rect 350552 16574 350580 177346
rect 350644 158710 350672 291178
rect 350724 252612 350776 252618
rect 350724 252554 350776 252560
rect 350632 158704 350684 158710
rect 350632 158646 350684 158652
rect 350736 153202 350764 252554
rect 350724 153196 350776 153202
rect 350724 153138 350776 153144
rect 351932 115938 351960 292538
rect 352024 142118 352052 295287
rect 352104 214600 352156 214606
rect 352104 214542 352156 214548
rect 352012 142112 352064 142118
rect 352012 142054 352064 142060
rect 351920 115932 351972 115938
rect 351920 115874 351972 115880
rect 352116 106282 352144 214542
rect 352104 106276 352156 106282
rect 352104 106218 352156 106224
rect 350552 16546 351224 16574
rect 350448 3528 350500 3534
rect 350448 3470 350500 3476
rect 350460 480 350488 3470
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 353312 3466 353340 389166
rect 395356 340202 395384 699654
rect 580262 683904 580318 683913
rect 580262 683839 580318 683848
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 580000 630698 580028 630799
rect 579988 630692 580040 630698
rect 579988 630634 580040 630640
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 579894 537840 579950 537849
rect 579894 537775 579950 537784
rect 579908 536858 579936 537775
rect 579896 536852 579948 536858
rect 579896 536794 579948 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580184 470626 580212 471407
rect 580172 470620 580224 470626
rect 580172 470562 580224 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 579894 431624 579950 431633
rect 579894 431559 579950 431568
rect 579908 430642 579936 431559
rect 579896 430636 579948 430642
rect 579896 430578 579948 430584
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580276 387122 580304 683839
rect 582378 617536 582434 617545
rect 582378 617471 582434 617480
rect 580264 387116 580316 387122
rect 580264 387058 580316 387064
rect 580262 378448 580318 378457
rect 580262 378383 580318 378392
rect 579618 365120 579674 365129
rect 579618 365055 579674 365064
rect 579632 364410 579660 365055
rect 579620 364404 579672 364410
rect 579620 364346 579672 364352
rect 580276 341562 580304 378383
rect 580356 362228 580408 362234
rect 580356 362170 580408 362176
rect 580368 351937 580396 362170
rect 580354 351928 580410 351937
rect 580354 351863 580410 351872
rect 580264 341556 580316 341562
rect 580264 341498 580316 341504
rect 395344 340196 395396 340202
rect 395344 340138 395396 340144
rect 582392 336054 582420 617471
rect 582380 336048 582432 336054
rect 582380 335990 582432 335996
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 317422 580212 325207
rect 582564 323604 582616 323610
rect 582564 323546 582616 323552
rect 580172 317416 580224 317422
rect 580172 317358 580224 317364
rect 580172 312588 580224 312594
rect 580172 312530 580224 312536
rect 580184 312089 580212 312530
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 356060 305040 356112 305046
rect 356060 304982 356112 304988
rect 353392 228404 353444 228410
rect 353392 228346 353444 228352
rect 353404 154562 353432 228346
rect 353392 154556 353444 154562
rect 353392 154498 353444 154504
rect 356072 121446 356100 304982
rect 582378 299568 582434 299577
rect 582378 299503 582434 299512
rect 580354 298752 580410 298761
rect 580354 298687 580410 298696
rect 358820 296744 358872 296750
rect 358820 296686 358872 296692
rect 357440 294024 357492 294030
rect 357440 293966 357492 293972
rect 356060 121440 356112 121446
rect 356060 121382 356112 121388
rect 357452 103494 357480 293966
rect 358832 122806 358860 296686
rect 580264 289128 580316 289134
rect 580264 289070 580316 289076
rect 468484 273964 468536 273970
rect 468484 273906 468536 273912
rect 464344 260160 464396 260166
rect 464344 260102 464396 260108
rect 464356 167006 464384 260102
rect 464344 167000 464396 167006
rect 464344 166942 464396 166948
rect 358820 122800 358872 122806
rect 358820 122742 358872 122748
rect 357440 103488 357492 103494
rect 357440 103430 357492 103436
rect 468496 100706 468524 273906
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 579896 259412 579948 259418
rect 579896 259354 579948 259360
rect 579908 258913 579936 259354
rect 579894 258904 579950 258913
rect 579894 258839 579950 258848
rect 580170 245576 580226 245585
rect 580170 245511 580226 245520
rect 580184 244322 580212 245511
rect 580172 244316 580224 244322
rect 580172 244258 580224 244264
rect 580276 179217 580304 289070
rect 580368 256018 580396 298687
rect 580540 269816 580592 269822
rect 580540 269758 580592 269764
rect 580448 265668 580500 265674
rect 580448 265610 580500 265616
rect 580356 256012 580408 256018
rect 580356 255954 580408 255960
rect 580356 247716 580408 247722
rect 580356 247658 580408 247664
rect 580262 179208 580318 179217
rect 580262 179143 580318 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580368 152697 580396 247658
rect 580460 205737 580488 265610
rect 580552 232393 580580 269758
rect 580538 232384 580594 232393
rect 580538 232319 580594 232328
rect 580446 205728 580502 205737
rect 580446 205663 580502 205672
rect 580354 152688 580410 152697
rect 580354 152623 580410 152632
rect 468484 100700 468536 100706
rect 468484 100642 468536 100648
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 582392 19825 582420 299503
rect 582470 298480 582526 298489
rect 582470 298415 582526 298424
rect 582484 73001 582512 298415
rect 582576 112849 582604 323546
rect 582840 308440 582892 308446
rect 582840 308382 582892 308388
rect 582748 233912 582800 233918
rect 582748 233854 582800 233860
rect 582656 195288 582708 195294
rect 582656 195230 582708 195236
rect 582562 112840 582618 112849
rect 582562 112775 582618 112784
rect 582470 72992 582526 73001
rect 582470 72927 582526 72936
rect 582378 19816 582434 19825
rect 582378 19751 582434 19760
rect 582668 6633 582696 195230
rect 582760 59673 582788 233854
rect 582852 219065 582880 308382
rect 583116 301504 583168 301510
rect 583116 301446 583168 301452
rect 582932 287700 582984 287706
rect 582932 287642 582984 287648
rect 582838 219056 582894 219065
rect 582838 218991 582894 219000
rect 582840 198008 582892 198014
rect 582840 197950 582892 197956
rect 582746 59664 582802 59673
rect 582746 59599 582802 59608
rect 582852 33153 582880 197950
rect 582944 126041 582972 287642
rect 583022 232520 583078 232529
rect 583022 232455 583078 232464
rect 582930 126032 582986 126041
rect 582930 125967 582986 125976
rect 583036 86193 583064 232455
rect 583128 192545 583156 301446
rect 583114 192536 583170 192545
rect 583114 192471 583170 192480
rect 583022 86184 583078 86193
rect 583022 86119 583078 86128
rect 582838 33144 582894 33153
rect 582838 33079 582894 33088
rect 582654 6624 582710 6633
rect 582654 6559 582710 6568
rect 353300 3460 353352 3466
rect 353300 3402 353352 3408
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632032 3478 632088
rect 3330 579944 3386 580000
rect 3238 566888 3294 566944
rect 2962 527856 3018 527912
rect 3054 501744 3110 501800
rect 3054 475632 3110 475688
rect 2778 462596 2834 462632
rect 2778 462576 2780 462596
rect 2780 462576 2832 462596
rect 2832 462576 2834 462596
rect 3146 449520 3202 449576
rect 2870 410488 2926 410544
rect 3330 371320 3386 371376
rect 3330 358400 3386 358456
rect 3330 345344 3386 345400
rect 3514 619112 3570 619168
rect 3514 606056 3570 606112
rect 3514 553852 3570 553888
rect 3514 553832 3516 553852
rect 3516 553832 3568 553852
rect 3568 553832 3570 553852
rect 3514 514820 3570 514856
rect 3514 514800 3516 514820
rect 3516 514800 3568 514820
rect 3568 514800 3570 514820
rect 3514 423544 3570 423600
rect 3514 397468 3516 397488
rect 3516 397468 3568 397488
rect 3568 397468 3570 397488
rect 3514 397432 3570 397468
rect 3514 319232 3570 319288
rect 3422 306176 3478 306232
rect 3330 267164 3386 267200
rect 3330 267144 3332 267164
rect 3332 267144 3384 267164
rect 3384 267144 3386 267164
rect 3146 254088 3202 254144
rect 3054 241032 3110 241088
rect 3330 214920 3386 214976
rect 1306 200640 1362 200696
rect 3238 162832 3294 162888
rect 2778 136720 2834 136776
rect 3146 110608 3202 110664
rect 3514 293120 3570 293176
rect 3606 201864 3662 201920
rect 3514 188808 3570 188864
rect 3514 149776 3570 149832
rect 3514 97552 3570 97608
rect 3514 84632 3570 84688
rect 3422 71576 3478 71632
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 2778 36488 2834 36544
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 4066 6432 4122 6488
rect 9678 12960 9734 13016
rect 22098 53080 22154 53136
rect 15198 4800 15254 4856
rect 49514 206216 49570 206272
rect 50986 238584 51042 238640
rect 52182 211792 52238 211848
rect 49698 62736 49754 62792
rect 53654 178608 53710 178664
rect 55034 238448 55090 238504
rect 57886 330384 57942 330440
rect 56598 64096 56654 64152
rect 60370 218592 60426 218648
rect 61658 253952 61714 254008
rect 61750 239400 61806 239456
rect 64694 297336 64750 297392
rect 60646 182824 60702 182880
rect 61934 93472 61990 93528
rect 67730 377032 67786 377088
rect 67638 376896 67694 376952
rect 67638 375672 67694 375728
rect 67546 375536 67602 375592
rect 67454 374312 67510 374368
rect 67362 374176 67418 374232
rect 66166 351872 66222 351928
rect 67638 373768 67694 373824
rect 67638 371728 67694 371784
rect 67638 368872 67694 368928
rect 67638 367512 67694 367568
rect 67638 365764 67694 365800
rect 67638 365744 67640 365764
rect 67640 365744 67692 365764
rect 67692 365744 67694 365764
rect 67730 364792 67786 364848
rect 67638 364420 67640 364440
rect 67640 364420 67692 364440
rect 67692 364420 67694 364440
rect 67638 364384 67694 364420
rect 67638 362072 67694 362128
rect 67638 360304 67694 360360
rect 67638 359352 67694 359408
rect 67730 359216 67786 359272
rect 67730 357992 67786 358048
rect 67638 357468 67694 357504
rect 67638 357448 67640 357468
rect 67640 357448 67692 357468
rect 67692 357448 67694 357468
rect 67638 356496 67694 356552
rect 67638 355272 67694 355328
rect 67730 354864 67786 354920
rect 67638 353912 67694 353968
rect 68098 353388 68154 353424
rect 68098 353368 68100 353388
rect 68100 353368 68152 353388
rect 68152 353368 68154 353388
rect 67638 352552 67694 352608
rect 68650 371864 68706 371920
rect 68558 363704 68614 363760
rect 68374 351872 68430 351928
rect 67638 351056 67694 351112
rect 67730 348472 67786 348528
rect 67638 348064 67694 348120
rect 67730 344664 67786 344720
rect 67638 344528 67694 344584
rect 67638 341672 67694 341728
rect 69110 369824 69166 369880
rect 69018 368464 69074 368520
rect 68834 363568 68890 363624
rect 68834 349152 68890 349208
rect 68742 342352 68798 342408
rect 68926 340176 68982 340232
rect 69202 349832 69258 349888
rect 72974 382336 73030 382392
rect 71686 379616 71742 379672
rect 74262 381112 74318 381168
rect 83278 381248 83334 381304
rect 89626 383696 89682 383752
rect 89810 380160 89866 380216
rect 94686 387776 94742 387832
rect 91742 383832 91798 383888
rect 91558 380976 91614 381032
rect 86958 379480 87014 379536
rect 71686 379380 71688 379400
rect 71688 379380 71740 379400
rect 71740 379380 71742 379400
rect 71686 379344 71742 379380
rect 108946 379344 109002 379400
rect 109498 379072 109554 379128
rect 109866 377712 109922 377768
rect 109774 373632 109830 373688
rect 110326 366560 110382 366616
rect 109590 360712 109646 360768
rect 109498 358128 109554 358184
rect 69294 345888 69350 345944
rect 70306 345888 70362 345944
rect 70490 340992 70546 341048
rect 69294 331880 69350 331936
rect 69202 325080 69258 325136
rect 67270 287952 67326 288008
rect 68742 293936 68798 293992
rect 68006 291080 68062 291136
rect 67546 290808 67602 290864
rect 67546 288496 67602 288552
rect 67454 287816 67510 287872
rect 67454 276256 67510 276312
rect 67730 287020 67786 287056
rect 67730 287000 67732 287020
rect 67732 287000 67784 287020
rect 67784 287000 67786 287020
rect 68190 285368 68246 285424
rect 70674 296792 70730 296848
rect 72422 313928 72478 313984
rect 71962 298288 72018 298344
rect 71042 292304 71098 292360
rect 73802 309712 73858 309768
rect 76562 339904 76618 339960
rect 75182 301416 75238 301472
rect 75182 295432 75238 295488
rect 75826 294072 75882 294128
rect 77390 337320 77446 337376
rect 77758 337320 77814 337376
rect 77114 293120 77170 293176
rect 82266 337456 82322 337512
rect 80978 335960 81034 336016
rect 81622 295296 81678 295352
rect 87602 324944 87658 325000
rect 88982 302776 89038 302832
rect 93214 304136 93270 304192
rect 91098 301552 91154 301608
rect 93950 300056 94006 300112
rect 90178 293256 90234 293312
rect 97722 334600 97778 334656
rect 102230 339360 102286 339416
rect 104162 333240 104218 333296
rect 105450 327664 105506 327720
rect 104806 305632 104862 305688
rect 106186 336640 106242 336696
rect 105818 299512 105874 299568
rect 110510 378120 110566 378176
rect 110418 358400 110474 358456
rect 110418 340720 110474 340776
rect 111798 378800 111854 378856
rect 111798 376796 111800 376816
rect 111800 376796 111852 376816
rect 111852 376796 111854 376816
rect 111798 376760 111854 376796
rect 111798 375400 111854 375456
rect 111798 374720 111854 374776
rect 111798 369980 111854 370016
rect 111798 369960 111800 369980
rect 111800 369960 111852 369980
rect 111852 369960 111854 369980
rect 111798 367240 111854 367296
rect 111798 365200 111854 365256
rect 110694 352960 110750 353016
rect 111062 352960 111118 353016
rect 110602 340720 110658 340776
rect 112074 376080 112130 376136
rect 111982 372680 112038 372736
rect 112442 373360 112498 373416
rect 112074 371320 112130 371376
rect 111982 367920 112038 367976
rect 111982 366288 112038 366344
rect 112350 372000 112406 372056
rect 113086 370640 113142 370696
rect 112166 365880 112222 365936
rect 111982 364520 112038 364576
rect 112074 363840 112130 363896
rect 111890 362480 111946 362536
rect 111982 361800 112038 361856
rect 111890 360440 111946 360496
rect 111982 359760 112038 359816
rect 111890 359080 111946 359136
rect 111890 357040 111946 357096
rect 111890 356360 111946 356416
rect 111890 355000 111946 355056
rect 111890 354320 111946 354376
rect 111890 351600 111946 351656
rect 111890 349560 111946 349616
rect 111890 348200 111946 348256
rect 111890 347520 111946 347576
rect 111890 345480 111946 345536
rect 111890 344800 111946 344856
rect 112074 355680 112130 355736
rect 111982 344120 112038 344176
rect 111890 343440 111946 343496
rect 111890 342080 111946 342136
rect 111890 340040 111946 340096
rect 112166 350240 112222 350296
rect 112258 348880 112314 348936
rect 113270 348880 113326 348936
rect 112166 346160 112222 346216
rect 113086 342760 113142 342816
rect 113178 340040 113234 340096
rect 114466 364928 114522 364984
rect 113822 357992 113878 358048
rect 113822 337320 113878 337376
rect 113822 319368 113878 319424
rect 113822 298424 113878 298480
rect 115294 382336 115350 382392
rect 115294 352552 115350 352608
rect 115294 294208 115350 294264
rect 114190 291896 114246 291952
rect 119986 343712 120042 343768
rect 116582 293392 116638 293448
rect 69018 291080 69074 291136
rect 68742 286048 68798 286104
rect 68650 284688 68706 284744
rect 68926 283736 68982 283792
rect 67638 283328 67694 283384
rect 67638 282104 67694 282160
rect 68282 280472 68338 280528
rect 67638 280336 67694 280392
rect 67730 279928 67786 279984
rect 67638 279248 67694 279304
rect 67730 277752 67786 277808
rect 67638 277616 67694 277672
rect 67638 276392 67694 276448
rect 67822 275032 67878 275088
rect 67638 274896 67694 274952
rect 67730 274488 67786 274544
rect 67822 272312 67878 272368
rect 67638 272176 67694 272232
rect 67638 270952 67694 271008
rect 67730 270816 67786 270872
rect 67730 269592 67786 269648
rect 67638 269456 67694 269512
rect 68190 268252 68246 268288
rect 68190 268232 68192 268252
rect 68192 268232 68244 268252
rect 68244 268232 68246 268252
rect 67638 268096 67694 268152
rect 67638 267588 67640 267608
rect 67640 267588 67692 267608
rect 67692 267588 67694 267608
rect 67638 267552 67694 267588
rect 67730 267008 67786 267064
rect 67730 265512 67786 265568
rect 67638 265376 67694 265432
rect 67638 264868 67640 264888
rect 67640 264868 67692 264888
rect 67692 264868 67694 264888
rect 67638 264832 67694 264868
rect 67730 263628 67786 263664
rect 67730 263608 67732 263628
rect 67732 263608 67784 263628
rect 67784 263608 67786 263628
rect 67638 263508 67640 263528
rect 67640 263508 67692 263528
rect 67692 263508 67694 263528
rect 67638 263472 67694 263508
rect 67638 262268 67694 262304
rect 67638 262248 67640 262268
rect 67640 262248 67692 262268
rect 67692 262248 67694 262268
rect 67638 261432 67694 261488
rect 67730 260908 67786 260944
rect 67730 260888 67732 260908
rect 67732 260888 67784 260908
rect 67784 260888 67786 260908
rect 67638 260788 67640 260808
rect 67640 260788 67692 260808
rect 67692 260788 67694 260808
rect 67638 260752 67694 260788
rect 67638 259528 67694 259584
rect 67730 258576 67786 258632
rect 67638 258188 67694 258224
rect 67638 258168 67640 258188
rect 67640 258168 67692 258188
rect 67692 258168 67694 258188
rect 67638 257896 67694 257952
rect 68374 273536 68430 273592
rect 67638 256808 67694 256864
rect 68834 255312 68890 255368
rect 67638 255212 67640 255232
rect 67640 255212 67692 255232
rect 67692 255212 67694 255232
rect 67638 255176 67694 255212
rect 67638 254496 67694 254552
rect 67638 253852 67640 253872
rect 67640 253852 67692 253872
rect 67692 253852 67694 253872
rect 67638 253816 67694 253852
rect 67638 252612 67694 252648
rect 67638 252592 67640 252612
rect 67640 252592 67692 252612
rect 67692 252592 67694 252612
rect 67730 251776 67786 251832
rect 67638 251252 67694 251288
rect 67638 251232 67640 251252
rect 67640 251232 67692 251252
rect 67692 251232 67694 251252
rect 67638 250416 67694 250472
rect 67730 249872 67786 249928
rect 67638 249756 67694 249792
rect 67638 249736 67640 249756
rect 67640 249736 67692 249756
rect 67692 249736 67694 249756
rect 68098 248668 68154 248704
rect 68098 248648 68100 248668
rect 68100 248648 68152 248668
rect 68152 248648 68154 248668
rect 67730 247696 67786 247752
rect 67638 247152 67694 247208
rect 67638 245248 67694 245304
rect 68098 244316 68154 244352
rect 68098 244296 68100 244316
rect 68100 244296 68152 244316
rect 68152 244296 68154 244316
rect 67638 243208 67694 243264
rect 67638 241848 67694 241904
rect 69018 255856 69074 255912
rect 120170 293256 120226 293312
rect 120170 285640 120226 285696
rect 120078 252320 120134 252376
rect 120078 250960 120134 251016
rect 120446 250996 120448 251016
rect 120448 250996 120500 251016
rect 120500 250996 120502 251016
rect 120446 250960 120502 250996
rect 69110 245656 69166 245712
rect 69202 243616 69258 243672
rect 69754 240216 69810 240272
rect 82082 239400 82138 239456
rect 86222 237224 86278 237280
rect 84382 226888 84438 226944
rect 91926 238448 91982 238504
rect 98366 238584 98422 238640
rect 74538 181328 74594 181384
rect 97262 179424 97318 179480
rect 99286 177656 99342 177712
rect 97262 176976 97318 177032
rect 104806 177656 104862 177712
rect 107566 177656 107622 177712
rect 110694 177656 110750 177712
rect 100666 176704 100722 176760
rect 102046 176724 102102 176760
rect 102046 176704 102048 176724
rect 102048 176704 102100 176724
rect 102100 176704 102102 176724
rect 103334 176704 103390 176760
rect 108118 176704 108174 176760
rect 110050 176704 110106 176760
rect 113822 238584 113878 238640
rect 117042 238448 117098 238504
rect 118962 239808 119018 239864
rect 121458 291760 121514 291816
rect 121458 291080 121514 291136
rect 121458 289756 121460 289776
rect 121460 289756 121512 289776
rect 121512 289756 121514 289776
rect 121458 289720 121514 289756
rect 121458 287680 121514 287736
rect 121458 287020 121514 287056
rect 121458 287000 121460 287020
rect 121460 287000 121512 287020
rect 121512 287000 121514 287020
rect 120814 285676 120816 285696
rect 120816 285676 120868 285696
rect 120868 285676 120870 285696
rect 120814 285640 120870 285676
rect 121550 286320 121606 286376
rect 121550 284960 121606 285016
rect 121458 283600 121514 283656
rect 121458 282940 121514 282976
rect 121458 282920 121460 282940
rect 121460 282920 121512 282940
rect 121512 282920 121514 282940
rect 121458 282240 121514 282296
rect 121550 280880 121606 280936
rect 121458 280236 121460 280256
rect 121460 280236 121512 280256
rect 121512 280236 121514 280256
rect 121458 280200 121514 280236
rect 121550 279520 121606 279576
rect 121458 278860 121514 278896
rect 121458 278840 121460 278860
rect 121460 278840 121512 278860
rect 121512 278840 121514 278860
rect 121550 278160 121606 278216
rect 121458 277500 121514 277536
rect 121458 277480 121460 277500
rect 121460 277480 121512 277500
rect 121512 277480 121514 277500
rect 121458 276800 121514 276856
rect 121458 276120 121514 276176
rect 121734 290400 121790 290456
rect 122286 289040 122342 289096
rect 121734 288360 121790 288416
rect 121734 284280 121790 284336
rect 121734 281560 121790 281616
rect 121642 275440 121698 275496
rect 121458 274080 121514 274136
rect 121458 273400 121514 273456
rect 121550 272720 121606 272776
rect 122102 272040 122158 272096
rect 121458 271360 121514 271416
rect 121642 270000 121698 270056
rect 121458 269320 121514 269376
rect 121550 268640 121606 268696
rect 121458 267960 121514 268016
rect 121550 267280 121606 267336
rect 121458 266600 121514 266656
rect 121550 265920 121606 265976
rect 121458 265240 121514 265296
rect 121458 264560 121514 264616
rect 121550 263880 121606 263936
rect 121458 263200 121514 263256
rect 121458 262520 121514 262576
rect 121550 261840 121606 261896
rect 121458 260480 121514 260536
rect 121458 259800 121514 259856
rect 121642 259120 121698 259176
rect 121550 258440 121606 258496
rect 121550 257760 121606 257816
rect 121458 257080 121514 257136
rect 121458 256400 121514 256456
rect 121550 255720 121606 255776
rect 121550 255040 121606 255096
rect 121458 254360 121514 254416
rect 121550 253680 121606 253736
rect 121458 253000 121514 253056
rect 121458 251640 121514 251696
rect 121550 250280 121606 250336
rect 121458 249600 121514 249656
rect 121550 248920 121606 248976
rect 121458 248240 121514 248296
rect 121642 247560 121698 247616
rect 121550 246880 121606 246936
rect 121458 246200 121514 246256
rect 121642 245520 121698 245576
rect 121550 244160 121606 244216
rect 121458 243480 121514 243536
rect 121734 244840 121790 244896
rect 121458 242836 121460 242856
rect 121460 242836 121512 242856
rect 121512 242836 121514 242856
rect 121458 242800 121514 242836
rect 121550 242120 121606 242176
rect 121458 240760 121514 240816
rect 121458 240080 121514 240136
rect 122746 261160 122802 261216
rect 124862 339360 124918 339416
rect 122930 241168 122986 241224
rect 125782 293392 125838 293448
rect 136730 351872 136786 351928
rect 140778 293120 140834 293176
rect 142802 351872 142858 351928
rect 114466 177656 114522 177712
rect 115846 177656 115902 177712
rect 116950 177656 117006 177712
rect 119986 177656 120042 177712
rect 120906 177656 120962 177712
rect 112166 176976 112222 177032
rect 125414 176976 125470 177032
rect 123298 176704 123354 176760
rect 159362 182960 159418 183016
rect 162122 379208 162178 379264
rect 129646 177656 129702 177712
rect 130750 177656 130806 177712
rect 166354 302776 166410 302832
rect 166354 179968 166410 180024
rect 162122 177248 162178 177304
rect 125874 176740 125876 176760
rect 125876 176740 125928 176760
rect 125928 176740 125930 176760
rect 125874 176704 125930 176740
rect 128266 176704 128322 176760
rect 133142 176704 133198 176760
rect 134430 176704 134486 176760
rect 136086 176704 136142 176760
rect 148230 176704 148286 176760
rect 127070 175480 127126 175536
rect 132038 175480 132094 175536
rect 158902 175480 158958 175536
rect 100758 175344 100814 175400
rect 118422 175344 118478 175400
rect 121918 175344 121974 175400
rect 167826 171536 167882 171592
rect 66166 129240 66222 129296
rect 65154 126248 65210 126304
rect 65522 125160 65578 125216
rect 66074 123528 66130 123584
rect 66074 102312 66130 102368
rect 67454 128016 67510 128072
rect 67362 122576 67418 122632
rect 66166 94832 66222 94888
rect 67546 120808 67602 120864
rect 67454 93744 67510 93800
rect 67638 100680 67694 100736
rect 129370 94696 129426 94752
rect 151726 94696 151782 94752
rect 85670 93608 85726 93664
rect 115478 93608 115534 93664
rect 120630 93608 120686 93664
rect 103426 93200 103482 93256
rect 110326 93200 110382 93256
rect 113822 93200 113878 93256
rect 74814 92420 74816 92440
rect 74816 92420 74868 92440
rect 74868 92420 74870 92440
rect 74814 92384 74870 92420
rect 88982 92404 89038 92440
rect 88982 92384 88984 92404
rect 88984 92384 89036 92404
rect 89036 92384 89038 92404
rect 95054 92384 95110 92440
rect 102046 92384 102102 92440
rect 99194 91296 99250 91352
rect 101862 91296 101918 91352
rect 85486 91160 85542 91216
rect 86866 91160 86922 91216
rect 88062 91160 88118 91216
rect 90730 91160 90786 91216
rect 92386 91160 92442 91216
rect 93766 91160 93822 91216
rect 95146 91160 95202 91216
rect 96526 91160 96582 91216
rect 97078 91160 97134 91216
rect 97906 91160 97962 91216
rect 66074 81368 66130 81424
rect 88062 86808 88118 86864
rect 99286 91160 99342 91216
rect 100206 91160 100262 91216
rect 100666 91160 100722 91216
rect 99286 80008 99342 80064
rect 101954 91160 102010 91216
rect 102966 91160 103022 91216
rect 105542 92384 105598 92440
rect 106646 92384 106702 92440
rect 106094 91704 106150 91760
rect 104806 91296 104862 91352
rect 104714 91160 104770 91216
rect 103426 84088 103482 84144
rect 77390 19896 77446 19952
rect 108210 91296 108266 91352
rect 109590 91296 109646 91352
rect 107198 91160 107254 91216
rect 106094 89664 106150 89720
rect 108486 91160 108542 91216
rect 110142 91160 110198 91216
rect 110694 91160 110750 91216
rect 111706 91160 111762 91216
rect 112534 91160 112590 91216
rect 110694 88168 110750 88224
rect 116766 92384 116822 92440
rect 135718 93608 135774 93664
rect 151726 93608 151782 93664
rect 128174 93200 128230 93256
rect 124034 92384 124090 92440
rect 115570 91704 115626 91760
rect 114466 91160 114522 91216
rect 122838 91432 122894 91488
rect 118238 91296 118294 91352
rect 119894 91296 119950 91352
rect 122654 91296 122710 91352
rect 115846 91160 115902 91216
rect 117134 91160 117190 91216
rect 118606 91160 118662 91216
rect 119986 91160 120042 91216
rect 121366 91160 121422 91216
rect 119894 83952 119950 84008
rect 122746 91160 122802 91216
rect 126702 92384 126758 92440
rect 134430 92384 134486 92440
rect 153014 92384 153070 92440
rect 126702 91976 126758 92032
rect 125414 91568 125470 91624
rect 124126 91160 124182 91216
rect 125506 91160 125562 91216
rect 126886 91568 126942 91624
rect 131026 91160 131082 91216
rect 132406 91160 132462 91216
rect 133234 91160 133290 91216
rect 151726 91160 151782 91216
rect 162858 89664 162914 89720
rect 168286 111732 168288 111752
rect 168288 111732 168340 111752
rect 168340 111732 168342 111752
rect 168286 111696 168342 111732
rect 167826 110064 167882 110120
rect 168102 108704 168158 108760
rect 178682 294072 178738 294128
rect 178682 95104 178738 95160
rect 178958 92248 179014 92304
rect 185582 177248 185638 177304
rect 189722 179968 189778 180024
rect 191194 182960 191250 183016
rect 195426 106800 195482 106856
rect 195334 93608 195390 93664
rect 199382 115096 199438 115152
rect 199566 93472 199622 93528
rect 210514 185544 210570 185600
rect 213918 176160 213974 176216
rect 213918 175072 213974 175128
rect 214010 174664 214066 174720
rect 213918 173712 213974 173768
rect 213918 172388 213920 172408
rect 213920 172388 213972 172408
rect 213972 172388 213974 172408
rect 213918 172352 213974 172388
rect 214010 171944 214066 172000
rect 214654 173304 214710 173360
rect 214470 170856 214526 170912
rect 213918 169652 213974 169688
rect 213918 169632 213920 169652
rect 213920 169632 213972 169652
rect 213972 169632 213974 169652
rect 214010 169360 214066 169416
rect 213918 168292 213974 168328
rect 213918 168272 213920 168292
rect 213920 168272 213972 168292
rect 213972 168272 213974 168292
rect 214010 168000 214066 168056
rect 214010 166640 214066 166696
rect 213918 166096 213974 166152
rect 213918 165280 213974 165336
rect 214010 164736 214066 164792
rect 213918 163376 213974 163432
rect 213918 162560 213974 162616
rect 214010 162016 214066 162072
rect 214930 170720 214986 170776
rect 214746 166912 214802 166968
rect 214654 161200 214710 161256
rect 213918 160792 213974 160848
rect 213918 158752 213974 158808
rect 213918 158652 213920 158672
rect 213920 158652 213972 158672
rect 213972 158652 213974 158672
rect 213918 158616 213974 158652
rect 214010 158072 214066 158128
rect 213918 157276 213974 157312
rect 213918 157256 213920 157276
rect 213920 157256 213972 157276
rect 213972 157256 213974 157276
rect 214010 156848 214066 156904
rect 213918 155916 213974 155952
rect 213918 155896 213920 155916
rect 213920 155896 213972 155916
rect 213972 155896 213974 155916
rect 214010 153856 214066 153912
rect 213918 153448 213974 153504
rect 214010 152632 214066 152688
rect 213918 151952 213974 152008
rect 214562 151816 214618 151872
rect 213918 150592 213974 150648
rect 214010 150048 214066 150104
rect 213918 148688 213974 148744
rect 213918 148008 213974 148064
rect 214010 146648 214066 146704
rect 213918 146376 213974 146432
rect 214010 145288 214066 145344
rect 213918 144880 213974 144936
rect 213918 143928 213974 143984
rect 214010 142704 214066 142760
rect 213918 142296 213974 142352
rect 213918 141344 213974 141400
rect 214010 140936 214066 140992
rect 214746 150728 214802 150784
rect 214654 149504 214710 149560
rect 214838 143520 214894 143576
rect 213274 139984 213330 140040
rect 213918 139460 213974 139496
rect 213918 139440 213920 139460
rect 213920 139440 213972 139460
rect 213972 139440 213974 139460
rect 213918 138080 213974 138136
rect 214470 137400 214526 137456
rect 213918 136720 213974 136776
rect 213918 135632 213974 135688
rect 213918 134000 213974 134056
rect 214010 132776 214066 132832
rect 213918 132524 213974 132560
rect 213918 132504 213920 132524
rect 213920 132504 213972 132524
rect 213972 132504 213974 132524
rect 214010 131416 214066 131472
rect 213918 131164 213974 131200
rect 213918 131144 213920 131164
rect 213920 131144 213972 131164
rect 213972 131144 213974 131164
rect 213918 129804 213974 129840
rect 213918 129784 213920 129804
rect 213920 129784 213972 129804
rect 213972 129784 213974 129804
rect 213918 128832 213974 128888
rect 213918 127064 213974 127120
rect 214010 126112 214066 126168
rect 213918 125724 213974 125760
rect 213918 125704 213920 125724
rect 213920 125704 213972 125724
rect 213972 125704 213974 125724
rect 214010 124752 214066 124808
rect 213918 124344 213974 124400
rect 214010 123528 214066 123584
rect 213918 123120 213974 123176
rect 214010 122168 214066 122224
rect 213918 121508 213974 121544
rect 213918 121488 213920 121508
rect 213920 121488 213972 121508
rect 213972 121488 213974 121508
rect 214010 120808 214066 120864
rect 213918 120400 213974 120456
rect 213366 119584 213422 119640
rect 214010 119040 214066 119096
rect 213918 118904 213974 118960
rect 214010 117544 214066 117600
rect 213918 117308 213920 117328
rect 213920 117308 213972 117328
rect 213972 117308 213974 117328
rect 213918 117272 213974 117308
rect 214010 116184 214066 116240
rect 213918 115948 213920 115968
rect 213920 115948 213972 115968
rect 213972 115948 213974 115968
rect 213918 115912 213974 115948
rect 213918 114960 213974 115016
rect 213918 113600 213974 113656
rect 213458 113192 213514 113248
rect 214010 112240 214066 112296
rect 213918 111852 213974 111888
rect 213918 111832 213920 111852
rect 213920 111832 213972 111852
rect 213972 111832 213974 111852
rect 214010 110880 214066 110936
rect 213918 110508 213920 110528
rect 213920 110508 213972 110528
rect 213972 110508 213974 110528
rect 213918 110472 213974 110508
rect 214010 109656 214066 109712
rect 213918 109248 213974 109304
rect 213918 107888 213974 107944
rect 214010 106936 214066 106992
rect 213918 106412 213974 106448
rect 213918 106392 213920 106412
rect 213920 106392 213972 106412
rect 213972 106392 213974 106412
rect 213918 105712 213974 105768
rect 214010 103944 214066 104000
rect 213918 103672 213974 103728
rect 214746 136040 214802 136096
rect 214654 108296 214710 108352
rect 215022 114552 215078 114608
rect 214010 102448 214066 102504
rect 213918 102312 213974 102368
rect 214010 101224 214066 101280
rect 213918 101088 213974 101144
rect 214102 99728 214158 99784
rect 214010 98368 214066 98424
rect 213918 97996 213920 98016
rect 213920 97996 213972 98016
rect 213972 97996 213974 98016
rect 213918 97960 213974 97996
rect 214562 96600 214618 96656
rect 214746 95784 214802 95840
rect 218702 192480 218758 192536
rect 229742 186904 229798 186960
rect 231122 177384 231178 177440
rect 232502 177248 232558 177304
rect 240782 178744 240838 178800
rect 240874 177520 240930 177576
rect 244922 176296 244978 176352
rect 242254 176160 242310 176216
rect 249246 175208 249302 175264
rect 249154 174256 249210 174312
rect 249154 172760 249210 172816
rect 249338 172352 249394 172408
rect 249798 166640 249854 166696
rect 250626 159296 250682 159352
rect 249890 153448 249946 153504
rect 249154 96600 249210 96656
rect 248418 26832 248474 26888
rect 252466 173712 252522 173768
rect 252466 171400 252522 171456
rect 251362 164328 251418 164384
rect 251270 159568 251326 159624
rect 252282 170448 252338 170504
rect 252466 170856 252522 170912
rect 252374 170040 252430 170096
rect 252466 169496 252522 169552
rect 252374 169088 252430 169144
rect 252466 168544 252522 168600
rect 252466 168136 252522 168192
rect 252466 167592 252522 167648
rect 252374 167184 252430 167240
rect 252466 166232 252522 166288
rect 252374 165688 252430 165744
rect 252466 165280 252522 165336
rect 252374 164736 252430 164792
rect 252374 163920 252430 163976
rect 252466 163376 252522 163432
rect 252282 162968 252338 163024
rect 252650 171808 252706 171864
rect 252558 162424 252614 162480
rect 252466 161472 252522 161528
rect 252466 161064 252522 161120
rect 252374 160520 252430 160576
rect 252006 160112 252062 160168
rect 252466 159160 252522 159216
rect 251454 158752 251510 158808
rect 252006 158616 252062 158672
rect 251178 157800 251234 157856
rect 251546 155352 251602 155408
rect 251362 150728 251418 150784
rect 251638 142704 251694 142760
rect 250626 136584 250682 136640
rect 251730 125704 251786 125760
rect 251822 115368 251878 115424
rect 252466 158208 252522 158264
rect 252466 156848 252522 156904
rect 252374 156304 252430 156360
rect 252466 155916 252522 155952
rect 252466 155896 252468 155916
rect 252468 155896 252520 155916
rect 252520 155896 252522 155916
rect 252466 154944 252522 155000
rect 252466 153992 252522 154048
rect 252466 153076 252468 153096
rect 252468 153076 252520 153096
rect 252520 153076 252522 153096
rect 252466 153040 252522 153076
rect 252374 152632 252430 152688
rect 252374 151700 252430 151736
rect 252374 151680 252376 151700
rect 252376 151680 252428 151700
rect 252428 151680 252430 151700
rect 252466 151136 252522 151192
rect 252098 149776 252154 149832
rect 252466 150184 252522 150240
rect 252282 149232 252338 149288
rect 252466 148824 252522 148880
rect 252374 148280 252430 148336
rect 252282 147872 252338 147928
rect 252834 154400 252890 154456
rect 252742 146920 252798 146976
rect 252466 146512 252522 146568
rect 252466 145968 252522 146024
rect 252374 145560 252430 145616
rect 252282 145016 252338 145072
rect 252190 144608 252246 144664
rect 252466 144064 252522 144120
rect 252374 143656 252430 143712
rect 252466 143112 252522 143168
rect 252374 142160 252430 142216
rect 253202 141616 253258 141672
rect 252466 141344 252522 141400
rect 252374 140800 252430 140856
rect 252006 140392 252062 140448
rect 252466 139848 252522 139904
rect 252374 139440 252430 139496
rect 252466 138896 252522 138952
rect 252374 138488 252430 138544
rect 252466 137536 252522 137592
rect 252374 136992 252430 137048
rect 252466 136176 252522 136232
rect 252374 135632 252430 135688
rect 252282 135224 252338 135280
rect 252466 134680 252522 134736
rect 252374 134272 252430 134328
rect 252466 133748 252522 133784
rect 252466 133728 252468 133748
rect 252468 133728 252520 133748
rect 252520 133728 252522 133748
rect 252374 133320 252430 133376
rect 252282 132776 252338 132832
rect 252466 132368 252522 132424
rect 252374 131824 252430 131880
rect 252282 131416 252338 131472
rect 252466 130872 252522 130928
rect 252374 130464 252430 130520
rect 252282 130056 252338 130112
rect 252098 129104 252154 129160
rect 252466 129512 252522 129568
rect 252374 128560 252430 128616
rect 252466 128152 252522 128208
rect 252282 127608 252338 127664
rect 252374 127200 252430 127256
rect 252466 126656 252522 126712
rect 252190 126248 252246 126304
rect 252282 125296 252338 125352
rect 252466 124752 252522 124808
rect 252374 124344 252430 124400
rect 252466 123936 252522 123992
rect 252374 123392 252430 123448
rect 252282 122984 252338 123040
rect 252466 122440 252522 122496
rect 252282 122032 252338 122088
rect 252374 121488 252430 121544
rect 252466 121080 252522 121136
rect 252374 120536 252430 120592
rect 252466 120128 252522 120184
rect 252466 119584 252522 119640
rect 252282 119176 252338 119232
rect 252006 118768 252062 118824
rect 252466 118224 252522 118280
rect 252466 117816 252522 117872
rect 252374 117272 252430 117328
rect 252466 116864 252522 116920
rect 252374 116320 252430 116376
rect 252466 115912 252522 115968
rect 252374 114960 252430 115016
rect 251914 114416 251970 114472
rect 251730 113464 251786 113520
rect 251730 108296 251786 108352
rect 251178 105984 251234 106040
rect 252466 114008 252522 114064
rect 252466 113092 252468 113112
rect 252468 113092 252520 113112
rect 252520 113092 252522 113112
rect 252466 113056 252522 113092
rect 252374 112648 252430 112704
rect 252466 112104 252522 112160
rect 252466 111732 252468 111752
rect 252468 111732 252520 111752
rect 252520 111732 252522 111752
rect 252466 111696 252522 111732
rect 252282 111152 252338 111208
rect 252374 110744 252430 110800
rect 252466 110200 252522 110256
rect 252374 109792 252430 109848
rect 252282 109248 252338 109304
rect 252466 108876 252468 108896
rect 252468 108876 252520 108896
rect 252520 108876 252522 108896
rect 252466 108840 252522 108876
rect 252374 107888 252430 107944
rect 252282 106936 252338 106992
rect 252466 107516 252468 107536
rect 252468 107516 252520 107536
rect 252520 107516 252522 107536
rect 252466 107480 252522 107516
rect 252374 106528 252430 106584
rect 252466 105576 252522 105632
rect 252190 105032 252246 105088
rect 252098 103672 252154 103728
rect 252190 102720 252246 102776
rect 252466 104080 252522 104136
rect 252466 103128 252522 103184
rect 252374 102176 252430 102232
rect 252282 101360 252338 101416
rect 252466 100816 252522 100872
rect 252466 100408 252522 100464
rect 252374 99864 252430 99920
rect 252282 99456 252338 99512
rect 253202 98912 253258 98968
rect 252466 98504 252522 98560
rect 252374 97960 252430 98016
rect 252190 97552 252246 97608
rect 251270 97008 251326 97064
rect 252466 97008 252522 97064
rect 251178 96192 251234 96248
rect 255318 80688 255374 80744
rect 251270 13096 251326 13152
rect 264518 131688 264574 131744
rect 258262 3440 258318 3496
rect 259458 3440 259514 3496
rect 264150 3440 264206 3496
rect 265346 3440 265402 3496
rect 266542 3440 266598 3496
rect 268842 3576 268898 3632
rect 273902 293120 273958 293176
rect 277122 3576 277178 3632
rect 279422 297336 279478 297392
rect 286598 3440 286654 3496
rect 290186 3576 290242 3632
rect 288990 3440 289046 3496
rect 295982 180104 296038 180160
rect 296074 175752 296130 175808
rect 296718 33768 296774 33824
rect 300214 179968 300270 180024
rect 307482 174800 307538 174856
rect 307574 174392 307630 174448
rect 307666 174020 307668 174040
rect 307668 174020 307720 174040
rect 307720 174020 307722 174040
rect 307666 173984 307722 174020
rect 307574 173576 307630 173632
rect 307482 173168 307538 173224
rect 307666 172624 307722 172680
rect 306562 172216 306618 172272
rect 307574 171808 307630 171864
rect 307666 171400 307722 171456
rect 307298 170992 307354 171048
rect 307666 170584 307722 170640
rect 307482 170176 307538 170232
rect 307390 169768 307446 169824
rect 307114 168408 307170 168464
rect 307298 168000 307354 168056
rect 307114 166368 307170 166424
rect 307022 165416 307078 165472
rect 305642 147736 305698 147792
rect 299478 14456 299534 14512
rect 299662 3304 299718 3360
rect 301962 3440 302018 3496
rect 303158 3440 303214 3496
rect 306746 163376 306802 163432
rect 306562 161200 306618 161256
rect 306930 158616 306986 158672
rect 306562 155624 306618 155680
rect 306562 154400 306618 154456
rect 306654 153176 306710 153232
rect 306562 152632 306618 152688
rect 306562 149776 306618 149832
rect 306930 146784 306986 146840
rect 306746 146376 306802 146432
rect 306562 144608 306618 144664
rect 306654 143792 306710 143848
rect 306470 142432 306526 142488
rect 306746 142704 306802 142760
rect 306654 141480 306710 141536
rect 307114 165008 307170 165064
rect 307574 169224 307630 169280
rect 307666 168816 307722 168872
rect 307482 167592 307538 167648
rect 307666 167184 307722 167240
rect 307574 166776 307630 166832
rect 307666 165824 307722 165880
rect 307206 164600 307262 164656
rect 307114 159568 307170 159624
rect 307666 164228 307668 164248
rect 307668 164228 307720 164248
rect 307720 164228 307722 164248
rect 307666 164192 307722 164228
rect 307574 163784 307630 163840
rect 307666 162968 307722 163024
rect 307482 162424 307538 162480
rect 307574 162016 307630 162072
rect 307666 161608 307722 161664
rect 307666 160792 307722 160848
rect 307574 160384 307630 160440
rect 307574 159976 307630 160032
rect 307666 159024 307722 159080
rect 307574 158208 307630 158264
rect 307390 157392 307446 157448
rect 307666 157800 307722 157856
rect 307482 156984 307538 157040
rect 307574 156576 307630 156632
rect 307666 156168 307722 156224
rect 307666 155216 307722 155272
rect 307206 154808 307262 154864
rect 307574 153992 307630 154048
rect 307666 153584 307722 153640
rect 307482 152224 307538 152280
rect 307666 151852 307668 151872
rect 307668 151852 307720 151872
rect 307720 151852 307722 151872
rect 307666 151816 307722 151852
rect 307482 151408 307538 151464
rect 307666 151000 307722 151056
rect 307574 150592 307630 150648
rect 307482 150184 307538 150240
rect 307574 149232 307630 149288
rect 307298 148824 307354 148880
rect 307390 147600 307446 147656
rect 307298 147192 307354 147248
rect 307666 148416 307722 148472
rect 307574 145832 307630 145888
rect 307482 145424 307538 145480
rect 307666 145016 307722 145072
rect 307666 144200 307722 144256
rect 307574 143384 307630 143440
rect 307666 142976 307722 143032
rect 307206 142024 307262 142080
rect 307114 141616 307170 141672
rect 306746 135632 306802 135688
rect 306562 133592 306618 133648
rect 307390 140800 307446 140856
rect 307298 139576 307354 139632
rect 307298 138216 307354 138272
rect 307206 136992 307262 137048
rect 306562 132232 306618 132288
rect 306930 131824 306986 131880
rect 306562 126792 306618 126848
rect 306562 125432 306618 125488
rect 306562 118632 306618 118688
rect 306930 116592 306986 116648
rect 307114 133184 307170 133240
rect 307114 121216 307170 121272
rect 307114 119992 307170 120048
rect 307114 117408 307170 117464
rect 307022 116184 307078 116240
rect 305826 108024 305882 108080
rect 305642 105304 305698 105360
rect 305734 101088 305790 101144
rect 306746 106800 306802 106856
rect 305918 106392 305974 106448
rect 306746 100000 306802 100056
rect 306930 97416 306986 97472
rect 306930 96192 306986 96248
rect 304354 3440 304410 3496
rect 305550 3440 305606 3496
rect 307114 115640 307170 115696
rect 307114 98640 307170 98696
rect 307666 140392 307722 140448
rect 307574 139032 307630 139088
rect 307666 138624 307722 138680
rect 307574 137808 307630 137864
rect 307666 137400 307722 137456
rect 307482 136584 307538 136640
rect 307574 136176 307630 136232
rect 307666 135224 307722 135280
rect 307666 134408 307722 134464
rect 307666 132640 307722 132696
rect 307482 131008 307538 131064
rect 307666 129920 307722 129976
rect 307298 129784 307354 129840
rect 307574 129240 307630 129296
rect 307482 128460 307484 128480
rect 307484 128460 307536 128480
rect 307536 128460 307538 128480
rect 307482 128424 307538 128460
rect 307666 128832 307722 128888
rect 307482 128016 307538 128072
rect 307574 127608 307630 127664
rect 307666 127200 307722 127256
rect 307666 125840 307722 125896
rect 307574 125024 307630 125080
rect 307482 124244 307484 124264
rect 307484 124244 307536 124264
rect 307536 124244 307538 124264
rect 307482 124208 307538 124244
rect 307666 124616 307722 124672
rect 307482 123800 307538 123856
rect 307574 123392 307630 123448
rect 307666 123004 307722 123040
rect 307666 122984 307668 123004
rect 307668 122984 307720 123004
rect 307720 122984 307722 123004
rect 307574 122440 307630 122496
rect 307482 121644 307538 121680
rect 307482 121624 307484 121644
rect 307484 121624 307536 121644
rect 307536 121624 307538 121644
rect 307666 122032 307722 122088
rect 307574 120808 307630 120864
rect 307666 120400 307722 120456
rect 307574 119584 307630 119640
rect 307666 119040 307722 119096
rect 307574 118224 307630 118280
rect 307666 117816 307722 117872
rect 307666 117000 307722 117056
rect 307574 115232 307630 115288
rect 307666 114824 307722 114880
rect 307482 114416 307538 114472
rect 307574 113600 307630 113656
rect 307666 113228 307668 113248
rect 307668 113228 307720 113248
rect 307720 113228 307722 113248
rect 307666 113192 307722 113228
rect 307666 112648 307722 112704
rect 307574 112240 307630 112296
rect 307666 111852 307722 111888
rect 307666 111832 307668 111852
rect 307668 111832 307720 111852
rect 307720 111832 307722 111852
rect 307574 111424 307630 111480
rect 307482 111016 307538 111072
rect 307666 110608 307722 110664
rect 307482 110200 307538 110256
rect 307574 109792 307630 109848
rect 307666 109248 307722 109304
rect 307666 108840 307722 108896
rect 307574 108432 307630 108488
rect 307482 107616 307538 107672
rect 307666 107208 307722 107264
rect 307574 105848 307630 105904
rect 307666 105052 307722 105088
rect 307666 105032 307668 105052
rect 307668 105032 307720 105052
rect 307720 105032 307722 105052
rect 307482 104624 307538 104680
rect 307574 104216 307630 104272
rect 307666 103808 307722 103864
rect 307482 103400 307538 103456
rect 307574 102992 307630 103048
rect 307666 102448 307722 102504
rect 307574 102040 307630 102096
rect 307482 100952 307538 101008
rect 307666 100852 307668 100872
rect 307668 100852 307720 100872
rect 307720 100852 307722 100872
rect 307666 100816 307722 100852
rect 307574 100408 307630 100464
rect 307666 99592 307722 99648
rect 307574 99048 307630 99104
rect 307666 98232 307722 98288
rect 307666 97824 307722 97880
rect 307666 96636 307668 96656
rect 307668 96636 307720 96656
rect 307720 96636 307722 96656
rect 307666 96600 307722 96636
rect 307850 30912 307906 30968
rect 308586 134816 308642 134872
rect 316682 253136 316738 253192
rect 313922 177384 313978 177440
rect 320822 175888 320878 175944
rect 321466 175208 321522 175264
rect 321282 169632 321338 169688
rect 321742 159840 321798 159896
rect 324594 217232 324650 217288
rect 321650 127472 321706 127528
rect 323030 181328 323086 181384
rect 324318 173984 324374 174040
rect 324318 173168 324374 173224
rect 324410 172352 324466 172408
rect 324318 170856 324374 170912
rect 323214 170040 323270 170096
rect 324318 168544 324374 168600
rect 324318 167728 324374 167784
rect 324410 167048 324466 167104
rect 324318 166232 324374 166288
rect 324318 165452 324320 165472
rect 324320 165452 324372 165472
rect 324372 165452 324374 165472
rect 324318 165416 324374 165452
rect 324410 164736 324466 164792
rect 324318 163920 324374 163976
rect 324410 163104 324466 163160
rect 324318 162424 324374 162480
rect 324410 161608 324466 161664
rect 324318 160792 324374 160848
rect 324410 160112 324466 160168
rect 324318 158480 324374 158536
rect 324410 157800 324466 157856
rect 324318 156984 324374 157040
rect 324318 156304 324374 156360
rect 324318 155488 324374 155544
rect 324410 154672 324466 154728
rect 324318 153992 324374 154048
rect 324318 153176 324374 153232
rect 324410 152360 324466 152416
rect 324318 151716 324320 151736
rect 324320 151716 324372 151736
rect 324372 151716 324374 151736
rect 324318 151680 324374 151716
rect 323122 150864 323178 150920
rect 324318 150048 324374 150104
rect 324410 149368 324466 149424
rect 324318 148552 324374 148608
rect 324318 147056 324374 147112
rect 324318 146260 324374 146296
rect 324318 146240 324320 146260
rect 324320 146240 324372 146260
rect 324372 146240 324374 146260
rect 324318 145424 324374 145480
rect 324318 144780 324320 144800
rect 324320 144780 324372 144800
rect 324372 144780 324374 144800
rect 324318 144744 324374 144780
rect 324410 143928 324466 143984
rect 324318 143112 324374 143168
rect 324410 142432 324466 142488
rect 324318 141616 324374 141672
rect 324318 140120 324374 140176
rect 324318 139340 324320 139360
rect 324320 139340 324372 139360
rect 324372 139340 324374 139360
rect 324318 139304 324374 139340
rect 324318 137844 324320 137864
rect 324320 137844 324372 137864
rect 324372 137844 324374 137864
rect 324318 137808 324374 137844
rect 324318 136348 324320 136368
rect 324320 136348 324372 136368
rect 324372 136348 324374 136368
rect 324318 136312 324374 136348
rect 324318 134680 324374 134736
rect 324318 133184 324374 133240
rect 324502 140800 324558 140856
rect 324502 138488 324558 138544
rect 324502 136992 324558 137048
rect 324502 135496 324558 135552
rect 324318 130872 324374 130928
rect 324410 130056 324466 130112
rect 324318 129376 324374 129432
rect 324410 128560 324466 128616
rect 324318 127744 324374 127800
rect 324502 126248 324558 126304
rect 324318 125432 324374 125488
rect 324318 123936 324374 123992
rect 324410 123120 324466 123176
rect 324318 122440 324374 122496
rect 323030 121624 323086 121680
rect 322938 120808 322994 120864
rect 324318 120128 324374 120184
rect 321558 119856 321614 119912
rect 324318 118532 324320 118552
rect 324320 118532 324372 118552
rect 324372 118532 324374 118552
rect 324318 118496 324374 118532
rect 324410 117816 324466 117872
rect 324318 116320 324374 116376
rect 324318 115504 324374 115560
rect 324410 114688 324466 114744
rect 324318 114008 324374 114064
rect 324410 113192 324466 113248
rect 324318 112376 324374 112432
rect 324318 110880 324374 110936
rect 324318 110064 324374 110120
rect 324410 109384 324466 109440
rect 324410 108568 324466 108624
rect 324318 107752 324374 107808
rect 324318 105440 324374 105496
rect 324318 104760 324374 104816
rect 324318 103164 324320 103184
rect 324320 103164 324372 103184
rect 324372 103164 324374 103184
rect 324318 103128 324374 103164
rect 321282 100408 321338 100464
rect 324318 100136 324374 100192
rect 321374 98776 321430 98832
rect 321558 97280 321614 97336
rect 321466 96600 321522 96656
rect 321374 95104 321430 95160
rect 324502 102448 324558 102504
rect 324962 132368 325018 132424
rect 325606 103944 325662 104000
rect 326066 175888 326122 175944
rect 326066 171128 326122 171184
rect 325882 147736 325938 147792
rect 324594 98504 324650 98560
rect 342258 298288 342314 298344
rect 319718 3440 319774 3496
rect 343822 182824 343878 182880
rect 346674 178608 346730 178664
rect 336278 3984 336334 4040
rect 335082 3576 335138 3632
rect 331586 3440 331642 3496
rect 332690 3440 332746 3496
rect 333886 3440 333942 3496
rect 337474 3440 337530 3496
rect 338670 3440 338726 3496
rect 339866 3440 339922 3496
rect 340970 3440 341026 3496
rect 343362 3440 343418 3496
rect 345754 3440 345810 3496
rect 352010 295296 352066 295352
rect 580262 683848 580318 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 579986 630808 580042 630864
rect 580170 590960 580226 591016
rect 580170 577632 580226 577688
rect 580170 564304 580226 564360
rect 579894 537784 579950 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 580170 471416 580226 471472
rect 580170 458088 580226 458144
rect 579894 431568 579950 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 582378 617480 582434 617536
rect 580262 378392 580318 378448
rect 579618 365064 579674 365120
rect 580354 351872 580410 351928
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 582378 299512 582434 299568
rect 580354 298696 580410 298752
rect 580170 272176 580226 272232
rect 579894 258848 579950 258904
rect 580170 245520 580226 245576
rect 580262 179152 580318 179208
rect 580170 165824 580226 165880
rect 580538 232328 580594 232384
rect 580446 205672 580502 205728
rect 580354 152632 580410 152688
rect 580170 99456 580226 99512
rect 580170 46280 580226 46336
rect 582470 298424 582526 298480
rect 582562 112784 582618 112840
rect 582470 72936 582526 72992
rect 582378 19760 582434 19816
rect 582838 219000 582894 219056
rect 582746 59608 582802 59664
rect 583022 232464 583078 232520
rect 582930 125976 582986 126032
rect 583114 192480 583170 192536
rect 583022 86128 583078 86184
rect 582838 33088 582894 33144
rect 582654 6568 582710 6624
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697234 584960 697324
rect 567150 697174 584960 697234
rect 69054 696900 69060 696964
rect 69124 696962 69130 696964
rect 567150 696962 567210 697174
rect 583520 697084 584960 697174
rect 69124 696902 567210 696962
rect 69124 696900 69130 696902
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580257 683906 580323 683909
rect 583520 683906 584960 683996
rect 580257 683904 584960 683906
rect 580257 683848 580262 683904
rect 580318 683848 584960 683904
rect 580257 683846 584960 683848
rect 580257 683843 580323 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 582373 617538 582439 617541
rect 583520 617538 584960 617628
rect 582373 617536 584960 617538
rect 582373 617480 582378 617536
rect 582434 617480 584960 617536
rect 582373 617478 584960 617480
rect 582373 617475 582439 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3233 566946 3299 566949
rect -960 566944 3299 566946
rect -960 566888 3238 566944
rect 3294 566888 3299 566944
rect -960 566886 3299 566888
rect -960 566796 480 566886
rect 3233 566883 3299 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3509 553890 3575 553893
rect -960 553888 3575 553890
rect -960 553832 3514 553888
rect 3570 553832 3575 553888
rect -960 553830 3575 553832
rect -960 553740 480 553830
rect 3509 553827 3575 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 579889 537842 579955 537845
rect 583520 537842 584960 537932
rect 579889 537840 584960 537842
rect 579889 537784 579894 537840
rect 579950 537784 584960 537840
rect 579889 537782 584960 537784
rect 579889 537779 579955 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3049 475690 3115 475693
rect -960 475688 3115 475690
rect -960 475632 3054 475688
rect 3110 475632 3115 475688
rect -960 475630 3115 475632
rect -960 475540 480 475630
rect 3049 475627 3115 475630
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 2773 462634 2839 462637
rect -960 462632 2839 462634
rect -960 462576 2778 462632
rect 2834 462576 2839 462632
rect -960 462574 2839 462576
rect -960 462484 480 462574
rect 2773 462571 2839 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 579889 431626 579955 431629
rect 583520 431626 584960 431716
rect 579889 431624 584960 431626
rect 579889 431568 579894 431624
rect 579950 431568 584960 431624
rect 579889 431566 584960 431568
rect 579889 431563 579955 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 2865 410546 2931 410549
rect -960 410544 2931 410546
rect -960 410488 2870 410544
rect 2926 410488 2931 410544
rect -960 410486 2931 410488
rect -960 410396 480 410486
rect 2865 410483 2931 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 583520 391628 584960 391868
rect 94681 387834 94747 387837
rect 177246 387834 177252 387836
rect 94681 387832 177252 387834
rect 94681 387776 94686 387832
rect 94742 387776 177252 387832
rect 94681 387774 177252 387776
rect 94681 387771 94747 387774
rect 177246 387772 177252 387774
rect 177316 387772 177322 387836
rect -960 384284 480 384524
rect 57830 383828 57836 383892
rect 57900 383890 57906 383892
rect 91737 383890 91803 383893
rect 57900 383888 91803 383890
rect 57900 383832 91742 383888
rect 91798 383832 91803 383888
rect 57900 383830 91803 383832
rect 57900 383828 57906 383830
rect 91737 383827 91803 383830
rect 89621 383754 89687 383757
rect 273846 383754 273852 383756
rect 89621 383752 273852 383754
rect 89621 383696 89626 383752
rect 89682 383696 273852 383752
rect 89621 383694 273852 383696
rect 89621 383691 89687 383694
rect 273846 383692 273852 383694
rect 273916 383692 273922 383756
rect 72969 382394 73035 382397
rect 115289 382394 115355 382397
rect 72969 382392 115355 382394
rect 72969 382336 72974 382392
rect 73030 382336 115294 382392
rect 115350 382336 115355 382392
rect 72969 382334 115355 382336
rect 72969 382331 73035 382334
rect 115289 382331 115355 382334
rect 83273 381306 83339 381309
rect 170254 381306 170260 381308
rect 83273 381304 170260 381306
rect 83273 381248 83278 381304
rect 83334 381248 170260 381304
rect 83273 381246 170260 381248
rect 83273 381243 83339 381246
rect 170254 381244 170260 381246
rect 170324 381244 170330 381308
rect 74257 381170 74323 381173
rect 262806 381170 262812 381172
rect 74257 381168 262812 381170
rect 74257 381112 74262 381168
rect 74318 381112 262812 381168
rect 74257 381110 262812 381112
rect 74257 381107 74323 381110
rect 262806 381108 262812 381110
rect 262876 381108 262882 381172
rect 91553 381034 91619 381037
rect 286174 381034 286180 381036
rect 91553 381032 286180 381034
rect 91553 380976 91558 381032
rect 91614 380976 286180 381032
rect 91553 380974 286180 380976
rect 91553 380971 91619 380974
rect 286174 380972 286180 380974
rect 286244 380972 286250 381036
rect 89805 380218 89871 380221
rect 303654 380218 303660 380220
rect 89805 380216 303660 380218
rect 89805 380160 89810 380216
rect 89866 380160 303660 380216
rect 89805 380158 303660 380160
rect 89805 380155 89871 380158
rect 303654 380156 303660 380158
rect 303724 380156 303730 380220
rect 71681 379674 71747 379677
rect 70718 379672 71747 379674
rect 70718 379616 71686 379672
rect 71742 379616 71747 379672
rect 70718 379614 71747 379616
rect 70718 379508 70778 379614
rect 71681 379611 71747 379614
rect 86953 379538 87019 379541
rect 298686 379538 298692 379540
rect 86953 379536 298692 379538
rect 86953 379480 86958 379536
rect 87014 379480 298692 379536
rect 86953 379478 298692 379480
rect 86953 379475 87019 379478
rect 298686 379476 298692 379478
rect 298756 379476 298762 379540
rect 71681 379402 71747 379405
rect 70902 379400 71747 379402
rect 70902 379344 71686 379400
rect 71742 379344 71747 379400
rect 70902 379342 71747 379344
rect 70902 379266 70962 379342
rect 71681 379339 71747 379342
rect 108941 379402 109007 379405
rect 108941 379400 113190 379402
rect 108941 379344 108946 379400
rect 109002 379344 113190 379400
rect 108941 379342 113190 379344
rect 108941 379339 109007 379342
rect 70718 379206 70962 379266
rect 113130 379266 113190 379342
rect 162117 379266 162183 379269
rect 113130 379264 162183 379266
rect 113130 379208 162122 379264
rect 162178 379208 162183 379264
rect 113130 379206 162183 379208
rect 70718 378828 70778 379206
rect 162117 379203 162183 379206
rect 109493 379130 109559 379133
rect 259494 379130 259500 379132
rect 109493 379128 259500 379130
rect 109493 379072 109498 379128
rect 109554 379072 259500 379128
rect 109493 379070 259500 379072
rect 109493 379067 109559 379070
rect 259494 379068 259500 379070
rect 259564 379068 259570 379132
rect 111793 378858 111859 378861
rect 109940 378856 111859 378858
rect 109940 378800 111798 378856
rect 111854 378800 111859 378856
rect 109940 378798 111859 378800
rect 111793 378795 111859 378798
rect 580257 378450 580323 378453
rect 583520 378450 584960 378540
rect 580257 378448 584960 378450
rect 580257 378392 580262 378448
rect 580318 378392 584960 378448
rect 580257 378390 584960 378392
rect 580257 378387 580323 378390
rect 583520 378300 584960 378390
rect 110505 378178 110571 378181
rect 109940 378176 110571 378178
rect 109940 378120 110510 378176
rect 110566 378120 110571 378176
rect 109940 378118 110571 378120
rect 110505 378115 110571 378118
rect 109861 377770 109927 377773
rect 304942 377770 304948 377772
rect 109861 377768 304948 377770
rect 109861 377712 109866 377768
rect 109922 377712 304948 377768
rect 109861 377710 304948 377712
rect 109861 377707 109927 377710
rect 304942 377708 304948 377710
rect 305012 377708 305018 377772
rect 67725 377090 67791 377093
rect 70166 377090 70226 377468
rect 109358 377092 109418 377468
rect 67725 377088 70226 377090
rect 67725 377032 67730 377088
rect 67786 377032 70226 377088
rect 67725 377030 70226 377032
rect 67725 377027 67791 377030
rect 109350 377028 109356 377092
rect 109420 377028 109426 377092
rect 67633 376954 67699 376957
rect 67633 376952 70226 376954
rect 67633 376896 67638 376952
rect 67694 376896 70226 376952
rect 67633 376894 70226 376896
rect 67633 376891 67699 376894
rect 70166 376788 70226 376894
rect 111793 376818 111859 376821
rect 109940 376816 111859 376818
rect 109940 376760 111798 376816
rect 111854 376760 111859 376816
rect 109940 376758 111859 376760
rect 111793 376755 111859 376758
rect 112069 376138 112135 376141
rect 109940 376136 112135 376138
rect 67633 375730 67699 375733
rect 70166 375730 70226 376108
rect 109940 376080 112074 376136
rect 112130 376080 112135 376136
rect 109940 376078 112135 376080
rect 112069 376075 112135 376078
rect 67633 375728 70226 375730
rect 67633 375672 67638 375728
rect 67694 375672 70226 375728
rect 67633 375670 70226 375672
rect 67633 375667 67699 375670
rect 67541 375594 67607 375597
rect 67541 375592 70226 375594
rect 67541 375536 67546 375592
rect 67602 375536 70226 375592
rect 67541 375534 70226 375536
rect 67541 375531 67607 375534
rect 70166 375428 70226 375534
rect 111793 375458 111859 375461
rect 109940 375456 111859 375458
rect 109940 375400 111798 375456
rect 111854 375400 111859 375456
rect 109940 375398 111859 375400
rect 111793 375395 111859 375398
rect 111793 374778 111859 374781
rect 109940 374776 111859 374778
rect 67449 374370 67515 374373
rect 70166 374370 70226 374748
rect 109940 374720 111798 374776
rect 111854 374720 111859 374776
rect 109940 374718 111859 374720
rect 111793 374715 111859 374718
rect 67449 374368 70226 374370
rect 67449 374312 67454 374368
rect 67510 374312 70226 374368
rect 67449 374310 70226 374312
rect 67449 374307 67515 374310
rect 67357 374234 67423 374237
rect 67357 374232 70226 374234
rect 67357 374176 67362 374232
rect 67418 374176 70226 374232
rect 67357 374174 70226 374176
rect 67357 374171 67423 374174
rect 70166 374068 70226 374174
rect 67633 373826 67699 373829
rect 67633 373824 70226 373826
rect 67633 373768 67638 373824
rect 67694 373768 70226 373824
rect 67633 373766 70226 373768
rect 67633 373763 67699 373766
rect 70166 373388 70226 373766
rect 109769 373690 109835 373693
rect 178534 373690 178540 373692
rect 109769 373688 178540 373690
rect 109769 373632 109774 373688
rect 109830 373632 178540 373688
rect 109769 373630 178540 373632
rect 109769 373627 109835 373630
rect 178534 373628 178540 373630
rect 178604 373628 178610 373692
rect 110638 373418 110644 373420
rect 109940 373358 110644 373418
rect 110638 373356 110644 373358
rect 110708 373418 110714 373420
rect 112437 373418 112503 373421
rect 110708 373416 112503 373418
rect 110708 373360 112442 373416
rect 112498 373360 112503 373416
rect 110708 373358 112503 373360
rect 110708 373356 110714 373358
rect 112437 373355 112503 373358
rect 111977 372738 112043 372741
rect 109940 372736 112043 372738
rect 109940 372680 111982 372736
rect 112038 372680 112043 372736
rect 109940 372678 112043 372680
rect 111977 372675 112043 372678
rect 112345 372058 112411 372061
rect 109940 372056 112411 372058
rect 68645 371922 68711 371925
rect 70166 371922 70226 372028
rect 109940 372000 112350 372056
rect 112406 372000 112411 372056
rect 109940 371998 112411 372000
rect 112345 371995 112411 371998
rect 68645 371920 70226 371922
rect 68645 371864 68650 371920
rect 68706 371864 70226 371920
rect 68645 371862 70226 371864
rect 68645 371859 68711 371862
rect 67633 371786 67699 371789
rect 67633 371784 70226 371786
rect 67633 371728 67638 371784
rect 67694 371728 70226 371784
rect 67633 371726 70226 371728
rect 67633 371723 67699 371726
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect 70166 371348 70226 371726
rect 112069 371378 112135 371381
rect 109940 371376 112135 371378
rect -960 371318 3391 371320
rect 109940 371320 112074 371376
rect 112130 371320 112135 371376
rect 109940 371318 112135 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 112069 371315 112135 371318
rect 113081 370698 113147 370701
rect 109940 370696 113147 370698
rect 65926 370228 65932 370292
rect 65996 370290 66002 370292
rect 70166 370290 70226 370668
rect 109940 370640 113086 370696
rect 113142 370640 113147 370696
rect 109940 370638 113147 370640
rect 113081 370635 113147 370638
rect 65996 370230 70226 370290
rect 65996 370228 66002 370230
rect 111793 370018 111859 370021
rect 109940 370016 111859 370018
rect 69105 369882 69171 369885
rect 70166 369882 70226 369988
rect 109940 369960 111798 370016
rect 111854 369960 111859 370016
rect 109940 369958 111859 369960
rect 111793 369955 111859 369958
rect 69105 369880 70226 369882
rect 69105 369824 69110 369880
rect 69166 369824 70226 369880
rect 69105 369822 70226 369824
rect 69105 369819 69171 369822
rect 67633 368930 67699 368933
rect 70166 368930 70226 369308
rect 67633 368928 70226 368930
rect 67633 368872 67638 368928
rect 67694 368872 70226 368928
rect 67633 368870 70226 368872
rect 67633 368867 67699 368870
rect 109910 368658 109970 369308
rect 69013 368522 69079 368525
rect 70166 368522 70226 368628
rect 109910 368598 113190 368658
rect 69013 368520 70226 368522
rect 69013 368464 69018 368520
rect 69074 368464 70226 368520
rect 69013 368462 70226 368464
rect 113130 368522 113190 368598
rect 269614 368522 269620 368524
rect 113130 368462 269620 368522
rect 69013 368459 69079 368462
rect 269614 368460 269620 368462
rect 269684 368460 269690 368524
rect 111977 367978 112043 367981
rect 109940 367976 112043 367978
rect 67633 367570 67699 367573
rect 70166 367570 70226 367948
rect 109940 367920 111982 367976
rect 112038 367920 112043 367976
rect 109940 367918 112043 367920
rect 111977 367915 112043 367918
rect 67633 367568 70226 367570
rect 67633 367512 67638 367568
rect 67694 367512 70226 367568
rect 67633 367510 70226 367512
rect 67633 367507 67699 367510
rect 111793 367298 111859 367301
rect 109940 367296 111859 367298
rect 109940 367240 111798 367296
rect 111854 367240 111859 367296
rect 109940 367238 111859 367240
rect 111793 367235 111859 367238
rect 110321 366618 110387 366621
rect 109940 366616 110387 366618
rect 66662 366148 66668 366212
rect 66732 366210 66738 366212
rect 70166 366210 70226 366588
rect 109940 366560 110326 366616
rect 110382 366560 110387 366616
rect 109940 366558 110387 366560
rect 110321 366555 110387 366558
rect 111977 366346 112043 366349
rect 335854 366346 335860 366348
rect 111977 366344 335860 366346
rect 111977 366288 111982 366344
rect 112038 366288 335860 366344
rect 111977 366286 335860 366288
rect 111977 366283 112043 366286
rect 335854 366284 335860 366286
rect 335924 366284 335930 366348
rect 66732 366150 70226 366210
rect 66732 366148 66738 366150
rect 112161 365938 112227 365941
rect 109940 365936 112227 365938
rect 67633 365802 67699 365805
rect 70166 365802 70226 365908
rect 109940 365880 112166 365936
rect 112222 365880 112227 365936
rect 109940 365878 112227 365880
rect 112161 365875 112227 365878
rect 67633 365800 70226 365802
rect 67633 365744 67638 365800
rect 67694 365744 70226 365800
rect 67633 365742 70226 365744
rect 67633 365739 67699 365742
rect 111793 365258 111859 365261
rect 109940 365256 111859 365258
rect 67725 364850 67791 364853
rect 70166 364850 70226 365228
rect 109940 365200 111798 365256
rect 111854 365200 111859 365256
rect 109940 365198 111859 365200
rect 111793 365195 111859 365198
rect 579613 365122 579679 365125
rect 583520 365122 584960 365212
rect 579613 365120 584960 365122
rect 579613 365064 579618 365120
rect 579674 365064 584960 365120
rect 579613 365062 584960 365064
rect 579613 365059 579679 365062
rect 114461 364986 114527 364989
rect 267774 364986 267780 364988
rect 114461 364984 267780 364986
rect 114461 364928 114466 364984
rect 114522 364928 267780 364984
rect 114461 364926 267780 364928
rect 114461 364923 114527 364926
rect 267774 364924 267780 364926
rect 267844 364924 267850 364988
rect 583520 364972 584960 365062
rect 67725 364848 70226 364850
rect 67725 364792 67730 364848
rect 67786 364792 70226 364848
rect 67725 364790 70226 364792
rect 67725 364787 67791 364790
rect 111977 364578 112043 364581
rect 109940 364576 112043 364578
rect 67633 364442 67699 364445
rect 70166 364442 70226 364548
rect 109940 364520 111982 364576
rect 112038 364520 112043 364576
rect 109940 364518 112043 364520
rect 111977 364515 112043 364518
rect 67633 364440 70226 364442
rect 67633 364384 67638 364440
rect 67694 364384 70226 364440
rect 67633 364382 70226 364384
rect 67633 364379 67699 364382
rect 112069 363898 112135 363901
rect 109940 363896 112135 363898
rect 68553 363762 68619 363765
rect 70166 363762 70226 363868
rect 109940 363840 112074 363896
rect 112130 363840 112135 363896
rect 109940 363838 112135 363840
rect 112069 363835 112135 363838
rect 68553 363760 70226 363762
rect 68553 363704 68558 363760
rect 68614 363704 70226 363760
rect 68553 363702 70226 363704
rect 68553 363699 68619 363702
rect 68829 363626 68895 363629
rect 68829 363624 70226 363626
rect 68829 363568 68834 363624
rect 68890 363568 70226 363624
rect 68829 363566 70226 363568
rect 68829 363563 68895 363566
rect 70166 363188 70226 363566
rect 111885 362538 111951 362541
rect 109940 362536 111951 362538
rect 67633 362130 67699 362133
rect 70166 362130 70226 362508
rect 109940 362480 111890 362536
rect 111946 362480 111951 362536
rect 109940 362478 111951 362480
rect 111885 362475 111951 362478
rect 67633 362128 70226 362130
rect 67633 362072 67638 362128
rect 67694 362072 70226 362128
rect 67633 362070 70226 362072
rect 67633 362067 67699 362070
rect 111977 361858 112043 361861
rect 109940 361856 112043 361858
rect 109940 361800 111982 361856
rect 112038 361800 112043 361856
rect 109940 361798 112043 361800
rect 111977 361795 112043 361798
rect 70166 360770 70226 361148
rect 64830 360710 70226 360770
rect 109542 360773 109602 361148
rect 109542 360768 109651 360773
rect 109542 360712 109590 360768
rect 109646 360712 109651 360768
rect 109542 360710 109651 360712
rect 64638 360300 64644 360364
rect 64708 360362 64714 360364
rect 64830 360362 64890 360710
rect 109585 360707 109651 360710
rect 111885 360498 111951 360501
rect 109940 360496 111951 360498
rect 64708 360302 64890 360362
rect 67633 360362 67699 360365
rect 70166 360362 70226 360468
rect 109940 360440 111890 360496
rect 111946 360440 111951 360496
rect 109940 360438 111951 360440
rect 111885 360435 111951 360438
rect 67633 360360 70226 360362
rect 67633 360304 67638 360360
rect 67694 360304 70226 360360
rect 67633 360302 70226 360304
rect 64708 360300 64714 360302
rect 67633 360299 67699 360302
rect 111977 359818 112043 359821
rect 109940 359816 112043 359818
rect 67633 359410 67699 359413
rect 70166 359410 70226 359788
rect 109940 359760 111982 359816
rect 112038 359760 112043 359816
rect 109940 359758 112043 359760
rect 111977 359755 112043 359758
rect 67633 359408 70226 359410
rect 67633 359352 67638 359408
rect 67694 359352 70226 359408
rect 67633 359350 70226 359352
rect 67633 359347 67699 359350
rect 67725 359274 67791 359277
rect 67725 359272 70226 359274
rect 67725 359216 67730 359272
rect 67786 359216 70226 359272
rect 67725 359214 70226 359216
rect 67725 359211 67791 359214
rect 70166 359108 70226 359214
rect 111885 359138 111951 359141
rect 109940 359136 111951 359138
rect 109940 359080 111890 359136
rect 111946 359080 111951 359136
rect 109940 359078 111951 359080
rect 111885 359075 111951 359078
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect 110413 358458 110479 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect 109940 358456 110479 358458
rect 109940 358428 110418 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 67725 358050 67791 358053
rect 70166 358050 70226 358428
rect 109910 358400 110418 358428
rect 110474 358400 110479 358456
rect 109910 358398 110479 358400
rect 109493 358186 109559 358189
rect 109910 358186 109970 358398
rect 110413 358395 110479 358398
rect 109493 358184 109970 358186
rect 109493 358128 109498 358184
rect 109554 358128 109970 358184
rect 109493 358126 109970 358128
rect 109493 358123 109559 358126
rect 67725 358048 70226 358050
rect 67725 357992 67730 358048
rect 67786 357992 70226 358048
rect 67725 357990 70226 357992
rect 113817 358050 113883 358053
rect 276238 358050 276244 358052
rect 113817 358048 276244 358050
rect 113817 357992 113822 358048
rect 113878 357992 276244 358048
rect 113817 357990 276244 357992
rect 67725 357987 67791 357990
rect 113817 357987 113883 357990
rect 276238 357988 276244 357990
rect 276308 357988 276314 358052
rect 67633 357506 67699 357509
rect 70166 357506 70226 357748
rect 67633 357504 70226 357506
rect 67633 357448 67638 357504
rect 67694 357448 70226 357504
rect 67633 357446 70226 357448
rect 67633 357443 67699 357446
rect 111885 357098 111951 357101
rect 109940 357096 111951 357098
rect 67633 356554 67699 356557
rect 70166 356554 70226 357068
rect 109940 357040 111890 357096
rect 111946 357040 111951 357096
rect 109940 357038 111951 357040
rect 111885 357035 111951 357038
rect 67633 356552 70226 356554
rect 67633 356496 67638 356552
rect 67694 356496 70226 356552
rect 67633 356494 70226 356496
rect 67633 356491 67699 356494
rect 111885 356418 111951 356421
rect 109940 356416 111951 356418
rect 109940 356360 111890 356416
rect 111946 356360 111951 356416
rect 109940 356358 111951 356360
rect 111885 356355 111951 356358
rect 112069 355738 112135 355741
rect 109940 355736 112135 355738
rect 67633 355330 67699 355333
rect 70166 355330 70226 355708
rect 109940 355680 112074 355736
rect 112130 355680 112135 355736
rect 109940 355678 112135 355680
rect 112069 355675 112135 355678
rect 67633 355328 70226 355330
rect 67633 355272 67638 355328
rect 67694 355272 70226 355328
rect 67633 355270 70226 355272
rect 67633 355267 67699 355270
rect 111885 355058 111951 355061
rect 109940 355056 111951 355058
rect 67725 354922 67791 354925
rect 70166 354922 70226 355028
rect 109940 355000 111890 355056
rect 111946 355000 111951 355056
rect 109940 354998 111951 355000
rect 111885 354995 111951 354998
rect 67725 354920 70226 354922
rect 67725 354864 67730 354920
rect 67786 354864 70226 354920
rect 67725 354862 70226 354864
rect 67725 354859 67791 354862
rect 111885 354378 111951 354381
rect 109940 354376 111951 354378
rect 67633 353970 67699 353973
rect 70166 353970 70226 354348
rect 109940 354320 111890 354376
rect 111946 354320 111951 354376
rect 109940 354318 111951 354320
rect 111885 354315 111951 354318
rect 67633 353968 70226 353970
rect 67633 353912 67638 353968
rect 67694 353912 70226 353968
rect 67633 353910 70226 353912
rect 67633 353907 67699 353910
rect 68093 353426 68159 353429
rect 70166 353426 70226 353668
rect 109910 353562 109970 353668
rect 271086 353562 271092 353564
rect 109910 353502 271092 353562
rect 271086 353500 271092 353502
rect 271156 353500 271162 353564
rect 68093 353424 70226 353426
rect 68093 353368 68098 353424
rect 68154 353368 70226 353424
rect 68093 353366 70226 353368
rect 68093 353363 68159 353366
rect 110689 353018 110755 353021
rect 111057 353018 111123 353021
rect 109940 353016 111123 353018
rect 67633 352610 67699 352613
rect 70166 352610 70226 352988
rect 109940 352960 110694 353016
rect 110750 352960 111062 353016
rect 111118 352960 111123 353016
rect 109940 352958 111123 352960
rect 110689 352955 110755 352958
rect 111057 352955 111123 352958
rect 67633 352608 70226 352610
rect 67633 352552 67638 352608
rect 67694 352552 70226 352608
rect 67633 352550 70226 352552
rect 115289 352610 115355 352613
rect 301814 352610 301820 352612
rect 115289 352608 301820 352610
rect 115289 352552 115294 352608
rect 115350 352552 301820 352608
rect 115289 352550 301820 352552
rect 67633 352547 67699 352550
rect 115289 352547 115355 352550
rect 301814 352548 301820 352550
rect 301884 352548 301890 352612
rect 66161 351930 66227 351933
rect 68369 351930 68435 351933
rect 70166 351930 70226 352308
rect 136725 351930 136791 351933
rect 142797 351930 142863 351933
rect 66161 351928 70226 351930
rect 66161 351872 66166 351928
rect 66222 351872 68374 351928
rect 68430 351872 70226 351928
rect 66161 351870 70226 351872
rect 113130 351928 142863 351930
rect 113130 351872 136730 351928
rect 136786 351872 142802 351928
rect 142858 351872 142863 351928
rect 113130 351870 142863 351872
rect 66161 351867 66227 351870
rect 68369 351867 68435 351870
rect 111885 351658 111951 351661
rect 109940 351656 111951 351658
rect 67633 351114 67699 351117
rect 70166 351114 70226 351628
rect 109940 351600 111890 351656
rect 111946 351600 111951 351656
rect 109940 351598 111951 351600
rect 111885 351595 111951 351598
rect 113130 351386 113190 351870
rect 136725 351867 136791 351870
rect 142797 351867 142863 351870
rect 580349 351930 580415 351933
rect 583520 351930 584960 352020
rect 580349 351928 584960 351930
rect 580349 351872 580354 351928
rect 580410 351872 584960 351928
rect 580349 351870 584960 351872
rect 580349 351867 580415 351870
rect 583520 351780 584960 351870
rect 67633 351112 70226 351114
rect 67633 351056 67638 351112
rect 67694 351056 70226 351112
rect 67633 351054 70226 351056
rect 109910 351326 113190 351386
rect 67633 351051 67699 351054
rect 109910 350948 109970 351326
rect 112161 350298 112227 350301
rect 109940 350296 112227 350298
rect 69197 349890 69263 349893
rect 70166 349890 70226 350268
rect 109940 350240 112166 350296
rect 112222 350240 112227 350296
rect 109940 350238 112227 350240
rect 112161 350235 112227 350238
rect 69197 349888 70226 349890
rect 69197 349832 69202 349888
rect 69258 349832 70226 349888
rect 69197 349830 70226 349832
rect 69197 349827 69263 349830
rect 111885 349618 111951 349621
rect 109940 349616 111951 349618
rect 68829 349210 68895 349213
rect 70166 349210 70226 349588
rect 109940 349560 111890 349616
rect 111946 349560 111951 349616
rect 109940 349558 111951 349560
rect 111885 349555 111951 349558
rect 68829 349208 70226 349210
rect 68829 349152 68834 349208
rect 68890 349152 70226 349208
rect 68829 349150 70226 349152
rect 68829 349147 68895 349150
rect 112253 348938 112319 348941
rect 113265 348938 113331 348941
rect 109940 348936 113331 348938
rect 67725 348530 67791 348533
rect 70166 348530 70226 348908
rect 109940 348880 112258 348936
rect 112314 348880 113270 348936
rect 113326 348880 113331 348936
rect 109940 348878 113331 348880
rect 112253 348875 112319 348878
rect 113265 348875 113331 348878
rect 67725 348528 70226 348530
rect 67725 348472 67730 348528
rect 67786 348472 70226 348528
rect 67725 348470 70226 348472
rect 67725 348467 67791 348470
rect 111885 348258 111951 348261
rect 109940 348256 111951 348258
rect 67633 348122 67699 348125
rect 70166 348122 70226 348228
rect 109940 348200 111890 348256
rect 111946 348200 111951 348256
rect 109940 348198 111951 348200
rect 111885 348195 111951 348198
rect 67633 348120 70226 348122
rect 67633 348064 67638 348120
rect 67694 348064 70226 348120
rect 67633 348062 70226 348064
rect 67633 348059 67699 348062
rect 111885 347578 111951 347581
rect 109940 347576 111951 347578
rect 66110 347108 66116 347172
rect 66180 347170 66186 347172
rect 70166 347170 70226 347548
rect 109940 347520 111890 347576
rect 111946 347520 111951 347576
rect 109940 347518 111951 347520
rect 111885 347515 111951 347518
rect 66180 347110 70226 347170
rect 66180 347108 66186 347110
rect 62982 346564 62988 346628
rect 63052 346626 63058 346628
rect 70166 346626 70226 346868
rect 63052 346566 70226 346626
rect 63052 346564 63058 346566
rect 112161 346218 112227 346221
rect 109940 346216 112227 346218
rect 70350 345949 70410 346188
rect 109940 346160 112166 346216
rect 112222 346160 112227 346216
rect 109940 346158 112227 346160
rect 112161 346155 112227 346158
rect 69289 345946 69355 345949
rect 70301 345946 70410 345949
rect 69289 345944 70410 345946
rect 69289 345888 69294 345944
rect 69350 345888 70306 345944
rect 70362 345888 70410 345944
rect 69289 345886 70410 345888
rect 69289 345883 69355 345886
rect 70301 345883 70367 345886
rect 111885 345538 111951 345541
rect 109940 345536 111951 345538
rect -960 345402 480 345492
rect 109940 345480 111890 345536
rect 111946 345480 111951 345536
rect 109940 345478 111951 345480
rect 111885 345475 111951 345478
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 111885 344858 111951 344861
rect 109940 344856 111951 344858
rect 67725 344722 67791 344725
rect 70166 344722 70226 344828
rect 109940 344800 111890 344856
rect 111946 344800 111951 344856
rect 109940 344798 111951 344800
rect 111885 344795 111951 344798
rect 67725 344720 70226 344722
rect 67725 344664 67730 344720
rect 67786 344664 70226 344720
rect 67725 344662 70226 344664
rect 67725 344659 67791 344662
rect 67633 344586 67699 344589
rect 67633 344584 70226 344586
rect 67633 344528 67638 344584
rect 67694 344528 70226 344584
rect 67633 344526 70226 344528
rect 67633 344523 67699 344526
rect 70166 344148 70226 344526
rect 111977 344178 112043 344181
rect 109940 344176 112043 344178
rect 109940 344120 111982 344176
rect 112038 344120 112043 344176
rect 109940 344118 112043 344120
rect 111977 344115 112043 344118
rect 119981 343770 120047 343773
rect 125726 343770 125732 343772
rect 119981 343768 125732 343770
rect 119981 343712 119986 343768
rect 120042 343712 125732 343768
rect 119981 343710 125732 343712
rect 119981 343707 120047 343710
rect 125726 343708 125732 343710
rect 125796 343708 125802 343772
rect 69054 343572 69060 343636
rect 69124 343634 69130 343636
rect 69124 343574 70410 343634
rect 69124 343572 69130 343574
rect 70350 343092 70410 343574
rect 111885 343498 111951 343501
rect 109940 343496 111951 343498
rect 109940 343440 111890 343496
rect 111946 343440 111951 343496
rect 109940 343438 111951 343440
rect 111885 343435 111951 343438
rect 70342 343028 70348 343092
rect 70412 343028 70418 343092
rect 113081 342818 113147 342821
rect 109940 342816 113147 342818
rect 68737 342410 68803 342413
rect 70166 342410 70226 342788
rect 109940 342760 113086 342816
rect 113142 342760 113147 342816
rect 109940 342758 113147 342760
rect 113081 342755 113147 342758
rect 68737 342408 70226 342410
rect 68737 342352 68742 342408
rect 68798 342352 70226 342408
rect 68737 342350 70226 342352
rect 68737 342347 68803 342350
rect 111885 342138 111951 342141
rect 109940 342136 111951 342138
rect 67633 341730 67699 341733
rect 70166 341730 70226 342108
rect 109940 342080 111890 342136
rect 111946 342080 111951 342136
rect 109940 342078 111951 342080
rect 111885 342075 111951 342078
rect 67633 341728 70226 341730
rect 67633 341672 67638 341728
rect 67694 341672 70226 341728
rect 67633 341670 70226 341672
rect 67633 341667 67699 341670
rect 70534 341053 70594 341428
rect 70485 341048 70594 341053
rect 70485 340992 70490 341048
rect 70546 340992 70594 341048
rect 70485 340990 70594 340992
rect 70485 340987 70551 340990
rect 110413 340778 110479 340781
rect 110597 340778 110663 340781
rect 109940 340776 110663 340778
rect 68921 340234 68987 340237
rect 70166 340234 70226 340748
rect 109940 340720 110418 340776
rect 110474 340720 110602 340776
rect 110658 340720 110663 340776
rect 109940 340718 110663 340720
rect 110413 340715 110479 340718
rect 110597 340715 110663 340718
rect 68921 340232 70226 340234
rect 68921 340176 68926 340232
rect 68982 340176 70226 340232
rect 68921 340174 70226 340176
rect 68921 340171 68987 340174
rect 111885 340098 111951 340101
rect 109940 340096 111951 340098
rect 109940 340040 111890 340096
rect 111946 340040 111951 340096
rect 109940 340038 111951 340040
rect 111885 340035 111951 340038
rect 113173 340098 113239 340101
rect 331254 340098 331260 340100
rect 113173 340096 331260 340098
rect 113173 340040 113178 340096
rect 113234 340040 331260 340096
rect 113173 340038 331260 340040
rect 113173 340035 113239 340038
rect 331254 340036 331260 340038
rect 331324 340036 331330 340100
rect 65926 339900 65932 339964
rect 65996 339962 66002 339964
rect 76557 339962 76623 339965
rect 65996 339960 76623 339962
rect 65996 339904 76562 339960
rect 76618 339904 76623 339960
rect 65996 339902 76623 339904
rect 65996 339900 66002 339902
rect 76557 339899 76623 339902
rect 102225 339418 102291 339421
rect 124254 339418 124260 339420
rect 102225 339416 124260 339418
rect 102225 339360 102230 339416
rect 102286 339360 124260 339416
rect 102225 339358 124260 339360
rect 102225 339355 102291 339358
rect 124254 339356 124260 339358
rect 124324 339418 124330 339420
rect 124857 339418 124923 339421
rect 124324 339416 124923 339418
rect 124324 339360 124862 339416
rect 124918 339360 124923 339416
rect 124324 339358 124923 339360
rect 124324 339356 124330 339358
rect 124857 339355 124923 339358
rect 583520 338452 584960 338692
rect 61878 337452 61884 337516
rect 61948 337514 61954 337516
rect 82261 337514 82327 337517
rect 61948 337512 82327 337514
rect 61948 337456 82266 337512
rect 82322 337456 82327 337512
rect 61948 337454 82327 337456
rect 61948 337452 61954 337454
rect 82261 337451 82327 337454
rect 70342 337316 70348 337380
rect 70412 337378 70418 337380
rect 77385 337378 77451 337381
rect 70412 337376 77451 337378
rect 70412 337320 77390 337376
rect 77446 337320 77451 337376
rect 70412 337318 77451 337320
rect 70412 337316 70418 337318
rect 77385 337315 77451 337318
rect 77753 337378 77819 337381
rect 113817 337378 113883 337381
rect 77753 337376 113883 337378
rect 77753 337320 77758 337376
rect 77814 337320 113822 337376
rect 113878 337320 113883 337376
rect 77753 337318 113883 337320
rect 77753 337315 77819 337318
rect 113817 337315 113883 337318
rect 106181 336698 106247 336701
rect 108982 336698 108988 336700
rect 106181 336696 108988 336698
rect 106181 336640 106186 336696
rect 106242 336640 108988 336696
rect 106181 336638 108988 336640
rect 106181 336635 106247 336638
rect 108982 336636 108988 336638
rect 109052 336636 109058 336700
rect 58934 335956 58940 336020
rect 59004 336018 59010 336020
rect 80973 336018 81039 336021
rect 59004 336016 81039 336018
rect 59004 335960 80978 336016
rect 81034 335960 81039 336016
rect 59004 335958 81039 335960
rect 59004 335956 59010 335958
rect 80973 335955 81039 335958
rect 97717 334658 97783 334661
rect 266302 334658 266308 334660
rect 97717 334656 266308 334658
rect 97717 334600 97722 334656
rect 97778 334600 266308 334656
rect 97717 334598 266308 334600
rect 97717 334595 97783 334598
rect 266302 334596 266308 334598
rect 266372 334596 266378 334660
rect 59118 333236 59124 333300
rect 59188 333298 59194 333300
rect 104157 333298 104223 333301
rect 59188 333296 104223 333298
rect 59188 333240 104162 333296
rect 104218 333240 104223 333296
rect 59188 333238 104223 333240
rect 59188 333236 59194 333238
rect 104157 333235 104223 333238
rect -960 332196 480 332436
rect 69289 331938 69355 331941
rect 118734 331938 118740 331940
rect 69289 331936 118740 331938
rect 69289 331880 69294 331936
rect 69350 331880 118740 331936
rect 69289 331878 118740 331880
rect 69289 331875 69355 331878
rect 118734 331876 118740 331878
rect 118804 331876 118810 331940
rect 66662 331740 66668 331804
rect 66732 331802 66738 331804
rect 338246 331802 338252 331804
rect 66732 331742 338252 331802
rect 66732 331740 66738 331742
rect 338246 331740 338252 331742
rect 338316 331740 338322 331804
rect 57881 330442 57947 330445
rect 263542 330442 263548 330444
rect 57881 330440 263548 330442
rect 57881 330384 57886 330440
rect 57942 330384 263548 330440
rect 57881 330382 263548 330384
rect 57881 330379 57947 330382
rect 263542 330380 263548 330382
rect 263612 330380 263618 330444
rect 105445 327722 105511 327725
rect 339534 327722 339540 327724
rect 105445 327720 339540 327722
rect 105445 327664 105450 327720
rect 105506 327664 339540 327720
rect 105445 327662 339540 327664
rect 105445 327659 105511 327662
rect 339534 327660 339540 327662
rect 339604 327660 339610 327724
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 69197 325138 69263 325141
rect 288382 325138 288388 325140
rect 69197 325136 288388 325138
rect 69197 325080 69202 325136
rect 69258 325080 288388 325136
rect 69197 325078 288388 325080
rect 69197 325075 69263 325078
rect 288382 325076 288388 325078
rect 288452 325076 288458 325140
rect 583520 325124 584960 325214
rect 87597 325002 87663 325005
rect 342294 325002 342300 325004
rect 87597 325000 342300 325002
rect 87597 324944 87602 325000
rect 87658 324944 342300 325000
rect 87597 324942 342300 324944
rect 87597 324939 87663 324942
rect 342294 324940 342300 324942
rect 342364 324940 342370 325004
rect 113817 319426 113883 319429
rect 340822 319426 340828 319428
rect 113817 319424 340828 319426
rect -960 319290 480 319380
rect 113817 319368 113822 319424
rect 113878 319368 340828 319424
rect 113817 319366 340828 319368
rect 113817 319363 113883 319366
rect 340822 319364 340828 319366
rect 340892 319364 340898 319428
rect 3509 319290 3575 319293
rect -960 319288 3575 319290
rect -960 319232 3514 319288
rect 3570 319232 3575 319288
rect -960 319230 3575 319232
rect -960 319140 480 319230
rect 3509 319227 3575 319230
rect 72417 313986 72483 313989
rect 265750 313986 265756 313988
rect 72417 313984 265756 313986
rect 72417 313928 72422 313984
rect 72478 313928 265756 313984
rect 72417 313926 265756 313928
rect 72417 313923 72483 313926
rect 265750 313924 265756 313926
rect 265820 313924 265826 313988
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect 73797 309770 73863 309773
rect 345054 309770 345060 309772
rect 73797 309768 345060 309770
rect 73797 309712 73802 309768
rect 73858 309712 345060 309768
rect 73797 309710 345060 309712
rect 73797 309707 73863 309710
rect 345054 309708 345060 309710
rect 345124 309708 345130 309772
rect -960 306234 480 306324
rect 3417 306234 3483 306237
rect -960 306232 3483 306234
rect -960 306176 3422 306232
rect 3478 306176 3483 306232
rect -960 306174 3483 306176
rect -960 306084 480 306174
rect 3417 306171 3483 306174
rect 104801 305690 104867 305693
rect 302182 305690 302188 305692
rect 104801 305688 302188 305690
rect 104801 305632 104806 305688
rect 104862 305632 302188 305688
rect 104801 305630 302188 305632
rect 104801 305627 104867 305630
rect 302182 305628 302188 305630
rect 302252 305628 302258 305692
rect 93209 304194 93275 304197
rect 334014 304194 334020 304196
rect 93209 304192 334020 304194
rect 93209 304136 93214 304192
rect 93270 304136 334020 304192
rect 93209 304134 334020 304136
rect 93209 304131 93275 304134
rect 334014 304132 334020 304134
rect 334084 304132 334090 304196
rect 88977 302834 89043 302837
rect 166349 302834 166415 302837
rect 88977 302832 166415 302834
rect 88977 302776 88982 302832
rect 89038 302776 166354 302832
rect 166410 302776 166415 302832
rect 88977 302774 166415 302776
rect 88977 302771 89043 302774
rect 166349 302771 166415 302774
rect 70894 301548 70900 301612
rect 70964 301610 70970 301612
rect 91093 301610 91159 301613
rect 70964 301608 91159 301610
rect 70964 301552 91098 301608
rect 91154 301552 91159 301608
rect 70964 301550 91159 301552
rect 70964 301548 70970 301550
rect 91093 301547 91159 301550
rect 75177 301474 75243 301477
rect 258390 301474 258396 301476
rect 75177 301472 258396 301474
rect 75177 301416 75182 301472
rect 75238 301416 258396 301472
rect 75177 301414 258396 301416
rect 75177 301411 75243 301414
rect 258390 301412 258396 301414
rect 258460 301412 258466 301476
rect 93945 300114 94011 300117
rect 110638 300114 110644 300116
rect 93945 300112 110644 300114
rect 93945 300056 93950 300112
rect 94006 300056 110644 300112
rect 93945 300054 110644 300056
rect 93945 300051 94011 300054
rect 110638 300052 110644 300054
rect 110708 300052 110714 300116
rect 105813 299570 105879 299573
rect 582373 299570 582439 299573
rect 105813 299568 582439 299570
rect 105813 299512 105818 299568
rect 105874 299512 582378 299568
rect 582434 299512 582439 299568
rect 105813 299510 582439 299512
rect 105813 299507 105879 299510
rect 582373 299507 582439 299510
rect 580349 298754 580415 298757
rect 583520 298754 584960 298844
rect 580349 298752 584960 298754
rect 580349 298696 580354 298752
rect 580410 298696 584960 298752
rect 580349 298694 584960 298696
rect 580349 298691 580415 298694
rect 583520 298604 584960 298694
rect 113817 298482 113883 298485
rect 582465 298482 582531 298485
rect 113817 298480 582531 298482
rect 113817 298424 113822 298480
rect 113878 298424 582470 298480
rect 582526 298424 582531 298480
rect 113817 298422 582531 298424
rect 113817 298419 113883 298422
rect 582465 298419 582531 298422
rect 71957 298346 72023 298349
rect 342253 298346 342319 298349
rect 71957 298344 342319 298346
rect 71957 298288 71962 298344
rect 72018 298288 342258 298344
rect 342314 298288 342319 298344
rect 71957 298286 342319 298288
rect 71957 298283 72023 298286
rect 342253 298283 342319 298286
rect 64689 297394 64755 297397
rect 279417 297394 279483 297397
rect 64689 297392 279483 297394
rect 64689 297336 64694 297392
rect 64750 297336 279422 297392
rect 279478 297336 279483 297392
rect 64689 297334 279483 297336
rect 64689 297331 64755 297334
rect 279417 297331 279483 297334
rect 70669 296850 70735 296853
rect 321502 296850 321508 296852
rect 70669 296848 321508 296850
rect 70669 296792 70674 296848
rect 70730 296792 321508 296848
rect 70669 296790 321508 296792
rect 70669 296787 70735 296790
rect 321502 296788 321508 296790
rect 321572 296788 321578 296852
rect 75177 295490 75243 295493
rect 252502 295490 252508 295492
rect 75177 295488 252508 295490
rect 75177 295432 75182 295488
rect 75238 295432 252508 295488
rect 75177 295430 252508 295432
rect 75177 295427 75243 295430
rect 252502 295428 252508 295430
rect 252572 295428 252578 295492
rect 81617 295354 81683 295357
rect 352005 295354 352071 295357
rect 81617 295352 352071 295354
rect 81617 295296 81622 295352
rect 81678 295296 352010 295352
rect 352066 295296 352071 295352
rect 81617 295294 352071 295296
rect 81617 295291 81683 295294
rect 352005 295291 352071 295294
rect 115289 294266 115355 294269
rect 123334 294266 123340 294268
rect 115289 294264 123340 294266
rect 115289 294208 115294 294264
rect 115350 294208 123340 294264
rect 115289 294206 123340 294208
rect 115289 294203 115355 294206
rect 123334 294204 123340 294206
rect 123404 294204 123410 294268
rect 75821 294130 75887 294133
rect 178677 294130 178743 294133
rect 75821 294128 178743 294130
rect 75821 294072 75826 294128
rect 75882 294072 178682 294128
rect 178738 294072 178743 294128
rect 75821 294070 178743 294072
rect 75821 294067 75887 294070
rect 178677 294067 178743 294070
rect 68737 293994 68803 293997
rect 322974 293994 322980 293996
rect 68737 293992 322980 293994
rect 68737 293936 68742 293992
rect 68798 293936 322980 293992
rect 68737 293934 322980 293936
rect 68737 293931 68803 293934
rect 322974 293932 322980 293934
rect 323044 293932 323050 293996
rect 116577 293450 116643 293453
rect 125777 293450 125843 293453
rect 116577 293448 125843 293450
rect 116577 293392 116582 293448
rect 116638 293392 125782 293448
rect 125838 293392 125843 293448
rect 116577 293390 125843 293392
rect 116577 293387 116643 293390
rect 125777 293387 125843 293390
rect 90173 293314 90239 293317
rect 120165 293314 120231 293317
rect 90173 293312 120231 293314
rect -960 293178 480 293268
rect 90173 293256 90178 293312
rect 90234 293256 120170 293312
rect 120226 293256 120231 293312
rect 90173 293254 120231 293256
rect 90173 293251 90239 293254
rect 120165 293251 120231 293254
rect 3509 293178 3575 293181
rect -960 293176 3575 293178
rect -960 293120 3514 293176
rect 3570 293120 3575 293176
rect -960 293118 3575 293120
rect -960 293028 480 293118
rect 3509 293115 3575 293118
rect 77109 293178 77175 293181
rect 140773 293178 140839 293181
rect 273897 293178 273963 293181
rect 77109 293176 273963 293178
rect 77109 293120 77114 293176
rect 77170 293120 140778 293176
rect 140834 293120 273902 293176
rect 273958 293120 273963 293176
rect 77109 293118 273963 293120
rect 77109 293115 77175 293118
rect 140773 293115 140839 293118
rect 273897 293115 273963 293118
rect 71037 292362 71103 292365
rect 70718 292360 71103 292362
rect 70718 292304 71042 292360
rect 71098 292304 71103 292360
rect 70718 292302 71103 292304
rect 70718 291788 70778 292302
rect 71037 292299 71103 292302
rect 114185 291954 114251 291957
rect 327022 291954 327028 291956
rect 114185 291952 327028 291954
rect 114185 291896 114190 291952
rect 114246 291896 327028 291952
rect 114185 291894 327028 291896
rect 114185 291891 114251 291894
rect 327022 291892 327028 291894
rect 327092 291892 327098 291956
rect 121453 291818 121519 291821
rect 119876 291816 121519 291818
rect 119876 291760 121458 291816
rect 121514 291760 121519 291816
rect 119876 291758 121519 291760
rect 121453 291755 121519 291758
rect 69982 291214 70226 291274
rect 68001 291138 68067 291141
rect 69013 291138 69079 291141
rect 69982 291138 70042 291214
rect 68001 291136 70042 291138
rect 68001 291080 68006 291136
rect 68062 291080 69018 291136
rect 69074 291080 70042 291136
rect 70166 291108 70226 291214
rect 121453 291138 121519 291141
rect 119876 291136 121519 291138
rect 68001 291078 70042 291080
rect 119876 291080 121458 291136
rect 121514 291080 121519 291136
rect 119876 291078 121519 291080
rect 68001 291075 68067 291078
rect 69013 291075 69079 291078
rect 121453 291075 121519 291078
rect 67541 290866 67607 290869
rect 67541 290864 70226 290866
rect 67541 290808 67546 290864
rect 67602 290808 70226 290864
rect 67541 290806 70226 290808
rect 67541 290803 67607 290806
rect 70166 290428 70226 290806
rect 121729 290458 121795 290461
rect 119876 290456 121795 290458
rect 119876 290400 121734 290456
rect 121790 290400 121795 290456
rect 119876 290398 121795 290400
rect 121729 290395 121795 290398
rect 121453 289778 121519 289781
rect 119876 289776 121519 289778
rect 65926 289172 65932 289236
rect 65996 289234 66002 289236
rect 70166 289234 70226 289748
rect 119876 289720 121458 289776
rect 121514 289720 121519 289776
rect 119876 289718 121519 289720
rect 121453 289715 121519 289718
rect 65996 289174 70226 289234
rect 65996 289172 66002 289174
rect 122281 289098 122347 289101
rect 119876 289096 122347 289098
rect 67541 288554 67607 288557
rect 70166 288554 70226 289068
rect 119876 289040 122286 289096
rect 122342 289040 122347 289096
rect 119876 289038 122347 289040
rect 122281 289035 122347 289038
rect 67541 288552 70226 288554
rect 67541 288496 67546 288552
rect 67602 288496 70226 288552
rect 67541 288494 70226 288496
rect 67541 288491 67607 288494
rect 121729 288418 121795 288421
rect 119876 288416 121795 288418
rect 67265 288010 67331 288013
rect 70350 288010 70410 288388
rect 119876 288360 121734 288416
rect 121790 288360 121795 288416
rect 119876 288358 121795 288360
rect 121729 288355 121795 288358
rect 67265 288008 70410 288010
rect 67265 287952 67270 288008
rect 67326 287952 70410 288008
rect 67265 287950 70410 287952
rect 67265 287947 67331 287950
rect 67449 287874 67515 287877
rect 67449 287872 70226 287874
rect 67449 287816 67454 287872
rect 67510 287816 70226 287872
rect 67449 287814 70226 287816
rect 67449 287811 67515 287814
rect 70166 287708 70226 287814
rect 121453 287738 121519 287741
rect 119876 287736 121519 287738
rect 119876 287680 121458 287736
rect 121514 287680 121519 287736
rect 119876 287678 121519 287680
rect 121453 287675 121519 287678
rect 67725 287058 67791 287061
rect 69982 287058 70226 287070
rect 121453 287058 121519 287061
rect 67725 287056 70226 287058
rect 67725 287000 67730 287056
rect 67786 287010 70226 287056
rect 119876 287056 121519 287058
rect 67786 287000 70042 287010
rect 67725 286998 70042 287000
rect 119876 287000 121458 287056
rect 121514 287000 121519 287056
rect 119876 286998 121519 287000
rect 67725 286995 67791 286998
rect 121453 286995 121519 286998
rect 70526 286724 70532 286788
rect 70596 286724 70602 286788
rect 70534 286348 70594 286724
rect 121545 286378 121611 286381
rect 119876 286376 121611 286378
rect 119876 286320 121550 286376
rect 121606 286320 121611 286376
rect 119876 286318 121611 286320
rect 121545 286315 121611 286318
rect 68737 286106 68803 286109
rect 68737 286104 70226 286106
rect 68737 286048 68742 286104
rect 68798 286048 70226 286104
rect 68737 286046 70226 286048
rect 68737 286043 68803 286046
rect 70166 285668 70226 286046
rect 120165 285698 120231 285701
rect 120809 285698 120875 285701
rect 119876 285696 120875 285698
rect 119876 285640 120170 285696
rect 120226 285640 120814 285696
rect 120870 285640 120875 285696
rect 119876 285638 120875 285640
rect 120165 285635 120231 285638
rect 120809 285635 120875 285638
rect 68185 285426 68251 285429
rect 68185 285424 70226 285426
rect 68185 285368 68190 285424
rect 68246 285368 70226 285424
rect 68185 285366 70226 285368
rect 68185 285363 68251 285366
rect 70166 284988 70226 285366
rect 583520 285276 584960 285516
rect 121545 285018 121611 285021
rect 119876 285016 121611 285018
rect 119876 284960 121550 285016
rect 121606 284960 121611 285016
rect 119876 284958 121611 284960
rect 121545 284955 121611 284958
rect 68645 284746 68711 284749
rect 68645 284744 70226 284746
rect 68645 284688 68650 284744
rect 68706 284688 70226 284744
rect 68645 284686 70226 284688
rect 68645 284683 68711 284686
rect 70166 284308 70226 284686
rect 121729 284338 121795 284341
rect 119876 284336 121795 284338
rect 119876 284280 121734 284336
rect 121790 284280 121795 284336
rect 119876 284278 121795 284280
rect 121729 284275 121795 284278
rect 68921 283794 68987 283797
rect 68921 283792 70226 283794
rect 68921 283736 68926 283792
rect 68982 283736 70226 283792
rect 68921 283734 70226 283736
rect 68921 283731 68987 283734
rect 70166 283628 70226 283734
rect 121453 283658 121519 283661
rect 119876 283656 121519 283658
rect 119876 283600 121458 283656
rect 121514 283600 121519 283656
rect 119876 283598 121519 283600
rect 121453 283595 121519 283598
rect 67633 283386 67699 283389
rect 67633 283384 70226 283386
rect 67633 283328 67638 283384
rect 67694 283328 70226 283384
rect 67633 283326 70226 283328
rect 67633 283323 67699 283326
rect 70166 282948 70226 283326
rect 121453 282978 121519 282981
rect 119876 282976 121519 282978
rect 119876 282920 121458 282976
rect 121514 282920 121519 282976
rect 119876 282918 121519 282920
rect 121453 282915 121519 282918
rect 121453 282298 121519 282301
rect 119876 282296 121519 282298
rect 119876 282240 121458 282296
rect 121514 282240 121519 282296
rect 119876 282238 121519 282240
rect 121453 282235 121519 282238
rect 67633 282162 67699 282165
rect 67633 282160 70226 282162
rect 67633 282104 67638 282160
rect 67694 282104 70226 282160
rect 67633 282102 70226 282104
rect 67633 282099 67699 282102
rect 70166 281588 70226 282102
rect 123334 282100 123340 282164
rect 123404 282162 123410 282164
rect 580206 282162 580212 282164
rect 123404 282102 580212 282162
rect 123404 282100 123410 282102
rect 580206 282100 580212 282102
rect 580276 282100 580282 282164
rect 121729 281618 121795 281621
rect 119876 281616 121795 281618
rect 119876 281560 121734 281616
rect 121790 281560 121795 281616
rect 119876 281558 121795 281560
rect 121729 281555 121795 281558
rect 121545 280938 121611 280941
rect 119876 280936 121611 280938
rect 68277 280530 68343 280533
rect 70166 280530 70226 280908
rect 119876 280880 121550 280936
rect 121606 280880 121611 280936
rect 119876 280878 121611 280880
rect 121545 280875 121611 280878
rect 68277 280528 70226 280530
rect 68277 280472 68282 280528
rect 68338 280472 70226 280528
rect 68277 280470 70226 280472
rect 68277 280467 68343 280470
rect 67633 280394 67699 280397
rect 67633 280392 70226 280394
rect 67633 280336 67638 280392
rect 67694 280336 70226 280392
rect 67633 280334 70226 280336
rect 67633 280331 67699 280334
rect 70166 280228 70226 280334
rect 121453 280258 121519 280261
rect 119876 280256 121519 280258
rect -960 279972 480 280212
rect 119876 280200 121458 280256
rect 121514 280200 121519 280256
rect 119876 280198 121519 280200
rect 121453 280195 121519 280198
rect 67725 279986 67791 279989
rect 67725 279984 70226 279986
rect 67725 279928 67730 279984
rect 67786 279928 70226 279984
rect 67725 279926 70226 279928
rect 67725 279923 67791 279926
rect 70166 279548 70226 279926
rect 121545 279578 121611 279581
rect 119876 279576 121611 279578
rect 119876 279520 121550 279576
rect 121606 279520 121611 279576
rect 119876 279518 121611 279520
rect 121545 279515 121611 279518
rect 67633 279306 67699 279309
rect 67633 279304 70226 279306
rect 67633 279248 67638 279304
rect 67694 279248 70226 279304
rect 67633 279246 70226 279248
rect 67633 279243 67699 279246
rect 70166 278868 70226 279246
rect 121453 278898 121519 278901
rect 119876 278896 121519 278898
rect 119876 278840 121458 278896
rect 121514 278840 121519 278896
rect 119876 278838 121519 278840
rect 121453 278835 121519 278838
rect 121545 278218 121611 278221
rect 119876 278216 121611 278218
rect 67725 277810 67791 277813
rect 70166 277810 70226 278188
rect 119876 278160 121550 278216
rect 121606 278160 121611 278216
rect 119876 278158 121611 278160
rect 121545 278155 121611 278158
rect 67725 277808 70226 277810
rect 67725 277752 67730 277808
rect 67786 277752 70226 277808
rect 67725 277750 70226 277752
rect 67725 277747 67791 277750
rect 67633 277674 67699 277677
rect 67633 277672 70226 277674
rect 67633 277616 67638 277672
rect 67694 277616 70226 277672
rect 67633 277614 70226 277616
rect 67633 277611 67699 277614
rect 70166 277508 70226 277614
rect 121453 277538 121519 277541
rect 119876 277536 121519 277538
rect 119876 277480 121458 277536
rect 121514 277480 121519 277536
rect 119876 277478 121519 277480
rect 121453 277475 121519 277478
rect 121453 276858 121519 276861
rect 119876 276856 121519 276858
rect 67633 276450 67699 276453
rect 70166 276450 70226 276828
rect 119876 276800 121458 276856
rect 121514 276800 121519 276856
rect 119876 276798 121519 276800
rect 121453 276795 121519 276798
rect 67633 276448 70226 276450
rect 67633 276392 67638 276448
rect 67694 276392 70226 276448
rect 67633 276390 70226 276392
rect 67633 276387 67699 276390
rect 67449 276314 67515 276317
rect 67449 276312 70226 276314
rect 67449 276256 67454 276312
rect 67510 276256 70226 276312
rect 67449 276254 70226 276256
rect 67449 276251 67515 276254
rect 70166 276148 70226 276254
rect 121453 276178 121519 276181
rect 119876 276176 121519 276178
rect 119876 276120 121458 276176
rect 121514 276120 121519 276176
rect 119876 276118 121519 276120
rect 121453 276115 121519 276118
rect 121637 275498 121703 275501
rect 119876 275496 121703 275498
rect 67817 275090 67883 275093
rect 70166 275090 70226 275468
rect 119876 275440 121642 275496
rect 121698 275440 121703 275496
rect 119876 275438 121703 275440
rect 121637 275435 121703 275438
rect 67817 275088 70226 275090
rect 67817 275032 67822 275088
rect 67878 275032 70226 275088
rect 67817 275030 70226 275032
rect 67817 275027 67883 275030
rect 67633 274954 67699 274957
rect 67633 274952 70226 274954
rect 67633 274896 67638 274952
rect 67694 274896 70226 274952
rect 67633 274894 70226 274896
rect 67633 274891 67699 274894
rect 70166 274788 70226 274894
rect 119876 274758 122850 274818
rect 122790 274682 122850 274758
rect 255262 274682 255268 274684
rect 122790 274622 255268 274682
rect 255262 274620 255268 274622
rect 255332 274620 255338 274684
rect 67725 274546 67791 274549
rect 67725 274544 70226 274546
rect 67725 274488 67730 274544
rect 67786 274488 70226 274544
rect 67725 274486 70226 274488
rect 67725 274483 67791 274486
rect 70166 274108 70226 274486
rect 121453 274138 121519 274141
rect 119876 274136 121519 274138
rect 119876 274080 121458 274136
rect 121514 274080 121519 274136
rect 119876 274078 121519 274080
rect 121453 274075 121519 274078
rect 68369 273594 68435 273597
rect 68369 273592 70226 273594
rect 68369 273536 68374 273592
rect 68430 273536 70226 273592
rect 68369 273534 70226 273536
rect 68369 273531 68435 273534
rect 70166 273428 70226 273534
rect 121453 273458 121519 273461
rect 119876 273456 121519 273458
rect 119876 273400 121458 273456
rect 121514 273400 121519 273456
rect 119876 273398 121519 273400
rect 121453 273395 121519 273398
rect 121545 272778 121611 272781
rect 119876 272776 121611 272778
rect 67817 272370 67883 272373
rect 70166 272370 70226 272748
rect 119876 272720 121550 272776
rect 121606 272720 121611 272776
rect 119876 272718 121611 272720
rect 121545 272715 121611 272718
rect 67817 272368 70226 272370
rect 67817 272312 67822 272368
rect 67878 272312 70226 272368
rect 67817 272310 70226 272312
rect 67817 272307 67883 272310
rect 67633 272234 67699 272237
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 67633 272232 70226 272234
rect 67633 272176 67638 272232
rect 67694 272176 70226 272232
rect 67633 272174 70226 272176
rect 67633 272171 67699 272174
rect 70166 272068 70226 272174
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 122097 272098 122163 272101
rect 119876 272096 122163 272098
rect 119876 272040 122102 272096
rect 122158 272040 122163 272096
rect 583520 272084 584960 272174
rect 119876 272038 122163 272040
rect 122097 272035 122163 272038
rect 121453 271418 121519 271421
rect 119876 271416 121519 271418
rect 67633 271010 67699 271013
rect 70166 271010 70226 271388
rect 119876 271360 121458 271416
rect 121514 271360 121519 271416
rect 119876 271358 121519 271360
rect 121453 271355 121519 271358
rect 67633 271008 70226 271010
rect 67633 270952 67638 271008
rect 67694 270952 70226 271008
rect 67633 270950 70226 270952
rect 67633 270947 67699 270950
rect 67725 270874 67791 270877
rect 67725 270872 70226 270874
rect 67725 270816 67730 270872
rect 67786 270816 70226 270872
rect 67725 270814 70226 270816
rect 67725 270811 67791 270814
rect 70166 270708 70226 270814
rect 121637 270058 121703 270061
rect 119876 270056 121703 270058
rect 67725 269650 67791 269653
rect 70166 269650 70226 270028
rect 119876 270000 121642 270056
rect 121698 270000 121703 270056
rect 119876 269998 121703 270000
rect 121637 269995 121703 269998
rect 67725 269648 70226 269650
rect 67725 269592 67730 269648
rect 67786 269592 70226 269648
rect 67725 269590 70226 269592
rect 67725 269587 67791 269590
rect 67633 269514 67699 269517
rect 67633 269512 70226 269514
rect 67633 269456 67638 269512
rect 67694 269456 70226 269512
rect 67633 269454 70226 269456
rect 67633 269451 67699 269454
rect 70166 269348 70226 269454
rect 121453 269378 121519 269381
rect 119876 269376 121519 269378
rect 119876 269320 121458 269376
rect 121514 269320 121519 269376
rect 119876 269318 121519 269320
rect 121453 269315 121519 269318
rect 121545 268698 121611 268701
rect 119876 268696 121611 268698
rect 68185 268290 68251 268293
rect 70166 268290 70226 268668
rect 119876 268640 121550 268696
rect 121606 268640 121611 268696
rect 119876 268638 121611 268640
rect 121545 268635 121611 268638
rect 68185 268288 70226 268290
rect 68185 268232 68190 268288
rect 68246 268232 70226 268288
rect 68185 268230 70226 268232
rect 68185 268227 68251 268230
rect 67633 268154 67699 268157
rect 67633 268152 70226 268154
rect 67633 268096 67638 268152
rect 67694 268096 70226 268152
rect 67633 268094 70226 268096
rect 67633 268091 67699 268094
rect 70166 267988 70226 268094
rect 121453 268018 121519 268021
rect 119876 268016 121519 268018
rect 119876 267960 121458 268016
rect 121514 267960 121519 268016
rect 119876 267958 121519 267960
rect 121453 267955 121519 267958
rect 67633 267610 67699 267613
rect 67633 267608 70226 267610
rect 67633 267552 67638 267608
rect 67694 267552 70226 267608
rect 67633 267550 70226 267552
rect 67633 267547 67699 267550
rect 70166 267308 70226 267550
rect 121545 267338 121611 267341
rect 119876 267336 121611 267338
rect -960 267202 480 267292
rect 119876 267280 121550 267336
rect 121606 267280 121611 267336
rect 119876 267278 121611 267280
rect 121545 267275 121611 267278
rect 3325 267202 3391 267205
rect -960 267200 3391 267202
rect -960 267144 3330 267200
rect 3386 267144 3391 267200
rect -960 267142 3391 267144
rect -960 267052 480 267142
rect 3325 267139 3391 267142
rect 67725 267066 67791 267069
rect 67725 267064 70226 267066
rect 67725 267008 67730 267064
rect 67786 267008 70226 267064
rect 67725 267006 70226 267008
rect 67725 267003 67791 267006
rect 70166 266628 70226 267006
rect 121453 266658 121519 266661
rect 119876 266656 121519 266658
rect 119876 266600 121458 266656
rect 121514 266600 121519 266656
rect 119876 266598 121519 266600
rect 121453 266595 121519 266598
rect 121545 265978 121611 265981
rect 119876 265976 121611 265978
rect 67725 265570 67791 265573
rect 70166 265570 70226 265948
rect 119876 265920 121550 265976
rect 121606 265920 121611 265976
rect 119876 265918 121611 265920
rect 121545 265915 121611 265918
rect 67725 265568 70226 265570
rect 67725 265512 67730 265568
rect 67786 265512 70226 265568
rect 67725 265510 70226 265512
rect 67725 265507 67791 265510
rect 67633 265434 67699 265437
rect 67633 265432 70226 265434
rect 67633 265376 67638 265432
rect 67694 265376 70226 265432
rect 67633 265374 70226 265376
rect 67633 265371 67699 265374
rect 70166 265268 70226 265374
rect 121453 265298 121519 265301
rect 119876 265296 121519 265298
rect 119876 265240 121458 265296
rect 121514 265240 121519 265296
rect 119876 265238 121519 265240
rect 121453 265235 121519 265238
rect 67633 264890 67699 264893
rect 67633 264888 70226 264890
rect 67633 264832 67638 264888
rect 67694 264832 70226 264888
rect 67633 264830 70226 264832
rect 67633 264827 67699 264830
rect 70166 264588 70226 264830
rect 121453 264618 121519 264621
rect 119876 264616 121519 264618
rect 119876 264560 121458 264616
rect 121514 264560 121519 264616
rect 119876 264558 121519 264560
rect 121453 264555 121519 264558
rect 121545 263938 121611 263941
rect 119876 263936 121611 263938
rect 67725 263666 67791 263669
rect 70166 263666 70226 263908
rect 119876 263880 121550 263936
rect 121606 263880 121611 263936
rect 119876 263878 121611 263880
rect 121545 263875 121611 263878
rect 67725 263664 70226 263666
rect 67725 263608 67730 263664
rect 67786 263608 70226 263664
rect 67725 263606 70226 263608
rect 67725 263603 67791 263606
rect 67633 263530 67699 263533
rect 67633 263528 70226 263530
rect 67633 263472 67638 263528
rect 67694 263472 70226 263528
rect 67633 263470 70226 263472
rect 67633 263467 67699 263470
rect 70166 263228 70226 263470
rect 121453 263258 121519 263261
rect 119876 263256 121519 263258
rect 119876 263200 121458 263256
rect 121514 263200 121519 263256
rect 119876 263198 121519 263200
rect 121453 263195 121519 263198
rect 121453 262578 121519 262581
rect 119876 262576 121519 262578
rect 67633 262306 67699 262309
rect 70166 262306 70226 262548
rect 119876 262520 121458 262576
rect 121514 262520 121519 262576
rect 119876 262518 121519 262520
rect 121453 262515 121519 262518
rect 67633 262304 70226 262306
rect 67633 262248 67638 262304
rect 67694 262248 70226 262304
rect 67633 262246 70226 262248
rect 67633 262243 67699 262246
rect 121545 261898 121611 261901
rect 119876 261896 121611 261898
rect 67633 261490 67699 261493
rect 70166 261490 70226 261868
rect 119876 261840 121550 261896
rect 121606 261840 121611 261896
rect 119876 261838 121611 261840
rect 121545 261835 121611 261838
rect 67633 261488 70226 261490
rect 67633 261432 67638 261488
rect 67694 261432 70226 261488
rect 67633 261430 70226 261432
rect 67633 261427 67699 261430
rect 122741 261218 122807 261221
rect 119876 261216 122807 261218
rect 67725 260946 67791 260949
rect 70166 260946 70226 261188
rect 119876 261160 122746 261216
rect 122802 261160 122807 261216
rect 119876 261158 122807 261160
rect 122741 261155 122807 261158
rect 67725 260944 70226 260946
rect 67725 260888 67730 260944
rect 67786 260888 70226 260944
rect 67725 260886 70226 260888
rect 67725 260883 67791 260886
rect 67633 260810 67699 260813
rect 67633 260808 70226 260810
rect 67633 260752 67638 260808
rect 67694 260752 70226 260808
rect 67633 260750 70226 260752
rect 67633 260747 67699 260750
rect 70166 260508 70226 260750
rect 121453 260538 121519 260541
rect 119876 260536 121519 260538
rect 119876 260480 121458 260536
rect 121514 260480 121519 260536
rect 119876 260478 121519 260480
rect 121453 260475 121519 260478
rect 121453 259858 121519 259861
rect 119876 259856 121519 259858
rect 67633 259586 67699 259589
rect 70350 259586 70410 259828
rect 119876 259800 121458 259856
rect 121514 259800 121519 259856
rect 119876 259798 121519 259800
rect 121453 259795 121519 259798
rect 67633 259584 70410 259586
rect 67633 259528 67638 259584
rect 67694 259528 70410 259584
rect 67633 259526 70410 259528
rect 67633 259523 67699 259526
rect 121637 259178 121703 259181
rect 119876 259176 121703 259178
rect 67725 258634 67791 258637
rect 70166 258634 70226 259148
rect 119876 259120 121642 259176
rect 121698 259120 121703 259176
rect 119876 259118 121703 259120
rect 121637 259115 121703 259118
rect 579889 258906 579955 258909
rect 583520 258906 584960 258996
rect 579889 258904 584960 258906
rect 579889 258848 579894 258904
rect 579950 258848 584960 258904
rect 579889 258846 584960 258848
rect 579889 258843 579955 258846
rect 583520 258756 584960 258846
rect 67725 258632 70226 258634
rect 67725 258576 67730 258632
rect 67786 258576 70226 258632
rect 67725 258574 70226 258576
rect 67725 258571 67791 258574
rect 121545 258498 121611 258501
rect 119876 258496 121611 258498
rect 67633 258226 67699 258229
rect 70166 258226 70226 258468
rect 119876 258440 121550 258496
rect 121606 258440 121611 258496
rect 119876 258438 121611 258440
rect 121545 258435 121611 258438
rect 67633 258224 70226 258226
rect 67633 258168 67638 258224
rect 67694 258168 70226 258224
rect 67633 258166 70226 258168
rect 67633 258163 67699 258166
rect 67633 257954 67699 257957
rect 67633 257952 70226 257954
rect 67633 257896 67638 257952
rect 67694 257896 70226 257952
rect 67633 257894 70226 257896
rect 67633 257891 67699 257894
rect 70166 257788 70226 257894
rect 121545 257818 121611 257821
rect 119876 257816 121611 257818
rect 119876 257760 121550 257816
rect 121606 257760 121611 257816
rect 119876 257758 121611 257760
rect 121545 257755 121611 257758
rect 121453 257138 121519 257141
rect 119876 257136 121519 257138
rect 67633 256866 67699 256869
rect 70350 256866 70410 257108
rect 119876 257080 121458 257136
rect 121514 257080 121519 257136
rect 119876 257078 121519 257080
rect 121453 257075 121519 257078
rect 67633 256864 70410 256866
rect 67633 256808 67638 256864
rect 67694 256808 70410 256864
rect 67633 256806 70410 256808
rect 67633 256803 67699 256806
rect 121453 256458 121519 256461
rect 119876 256456 121519 256458
rect 69013 255914 69079 255917
rect 70166 255914 70226 256428
rect 119876 256400 121458 256456
rect 121514 256400 121519 256456
rect 119876 256398 121519 256400
rect 121453 256395 121519 256398
rect 69013 255912 70226 255914
rect 69013 255856 69018 255912
rect 69074 255856 70226 255912
rect 69013 255854 70226 255856
rect 69013 255851 69079 255854
rect 121545 255778 121611 255781
rect 119876 255776 121611 255778
rect 68829 255370 68895 255373
rect 70166 255370 70226 255748
rect 119876 255720 121550 255776
rect 121606 255720 121611 255776
rect 119876 255718 121611 255720
rect 121545 255715 121611 255718
rect 68829 255368 70226 255370
rect 68829 255312 68834 255368
rect 68890 255312 70226 255368
rect 68829 255310 70226 255312
rect 68829 255307 68895 255310
rect 67633 255234 67699 255237
rect 67633 255232 70226 255234
rect 67633 255176 67638 255232
rect 67694 255176 70226 255232
rect 67633 255174 70226 255176
rect 67633 255171 67699 255174
rect 70166 255068 70226 255174
rect 121545 255098 121611 255101
rect 119876 255096 121611 255098
rect 119876 255040 121550 255096
rect 121606 255040 121611 255096
rect 119876 255038 121611 255040
rect 121545 255035 121611 255038
rect 67633 254554 67699 254557
rect 67633 254552 70226 254554
rect 67633 254496 67638 254552
rect 67694 254496 70226 254552
rect 67633 254494 70226 254496
rect 67633 254491 67699 254494
rect 70166 254388 70226 254494
rect 121453 254418 121519 254421
rect 119876 254416 121519 254418
rect 119876 254360 121458 254416
rect 121514 254360 121519 254416
rect 119876 254358 121519 254360
rect 121453 254355 121519 254358
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 61653 254012 61719 254013
rect 61653 254008 61700 254012
rect 61764 254010 61770 254012
rect 61653 253952 61658 254008
rect 61653 253948 61700 253952
rect 61764 253950 61810 254010
rect 61764 253948 61770 253950
rect 61653 253947 61719 253948
rect 67633 253874 67699 253877
rect 67633 253872 70226 253874
rect 67633 253816 67638 253872
rect 67694 253816 70226 253872
rect 67633 253814 70226 253816
rect 67633 253811 67699 253814
rect 70166 253708 70226 253814
rect 121545 253738 121611 253741
rect 119876 253736 121611 253738
rect 119876 253680 121550 253736
rect 121606 253680 121611 253736
rect 119876 253678 121611 253680
rect 121545 253675 121611 253678
rect 316677 253194 316743 253197
rect 332542 253194 332548 253196
rect 316677 253192 332548 253194
rect 316677 253136 316682 253192
rect 316738 253136 332548 253192
rect 316677 253134 332548 253136
rect 316677 253131 316743 253134
rect 332542 253132 332548 253134
rect 332612 253132 332618 253196
rect 121453 253058 121519 253061
rect 119876 253056 121519 253058
rect 67633 252650 67699 252653
rect 70166 252650 70226 253028
rect 119876 253000 121458 253056
rect 121514 253000 121519 253056
rect 119876 252998 121519 253000
rect 121453 252995 121519 252998
rect 67633 252648 70226 252650
rect 67633 252592 67638 252648
rect 67694 252592 70226 252648
rect 67633 252590 70226 252592
rect 67633 252587 67699 252590
rect 120073 252378 120139 252381
rect 119876 252376 120139 252378
rect 67725 251834 67791 251837
rect 70166 251834 70226 252348
rect 119876 252320 120078 252376
rect 120134 252320 120139 252376
rect 119876 252318 120139 252320
rect 120073 252315 120139 252318
rect 67725 251832 70226 251834
rect 67725 251776 67730 251832
rect 67786 251776 70226 251832
rect 67725 251774 70226 251776
rect 67725 251771 67791 251774
rect 121453 251698 121519 251701
rect 119876 251696 121519 251698
rect 67633 251290 67699 251293
rect 70166 251290 70226 251668
rect 119876 251640 121458 251696
rect 121514 251640 121519 251696
rect 119876 251638 121519 251640
rect 121453 251635 121519 251638
rect 67633 251288 70226 251290
rect 67633 251232 67638 251288
rect 67694 251232 70226 251288
rect 67633 251230 70226 251232
rect 67633 251227 67699 251230
rect 120073 251018 120139 251021
rect 120441 251018 120507 251021
rect 119876 251016 120507 251018
rect 67633 250474 67699 250477
rect 70166 250474 70226 250988
rect 119876 250960 120078 251016
rect 120134 250960 120446 251016
rect 120502 250960 120507 251016
rect 119876 250958 120507 250960
rect 120073 250955 120139 250958
rect 120441 250955 120507 250958
rect 67633 250472 70226 250474
rect 67633 250416 67638 250472
rect 67694 250416 70226 250472
rect 67633 250414 70226 250416
rect 67633 250411 67699 250414
rect 121545 250338 121611 250341
rect 119876 250336 121611 250338
rect 67725 249930 67791 249933
rect 70166 249930 70226 250308
rect 119876 250280 121550 250336
rect 121606 250280 121611 250336
rect 119876 250278 121611 250280
rect 121545 250275 121611 250278
rect 67725 249928 70226 249930
rect 67725 249872 67730 249928
rect 67786 249872 70226 249928
rect 67725 249870 70226 249872
rect 67725 249867 67791 249870
rect 67633 249794 67699 249797
rect 67633 249792 70226 249794
rect 67633 249736 67638 249792
rect 67694 249736 70226 249792
rect 67633 249734 70226 249736
rect 67633 249731 67699 249734
rect 70166 249628 70226 249734
rect 121453 249658 121519 249661
rect 119876 249656 121519 249658
rect 119876 249600 121458 249656
rect 121514 249600 121519 249656
rect 119876 249598 121519 249600
rect 121453 249595 121519 249598
rect 121545 248978 121611 248981
rect 119876 248976 121611 248978
rect 68093 248706 68159 248709
rect 70166 248706 70226 248948
rect 119876 248920 121550 248976
rect 121606 248920 121611 248976
rect 119876 248918 121611 248920
rect 121545 248915 121611 248918
rect 68093 248704 70226 248706
rect 68093 248648 68098 248704
rect 68154 248648 70226 248704
rect 68093 248646 70226 248648
rect 68093 248643 68159 248646
rect 121453 248298 121519 248301
rect 119876 248296 121519 248298
rect 67725 247754 67791 247757
rect 70166 247754 70226 248268
rect 119876 248240 121458 248296
rect 121514 248240 121519 248296
rect 119876 248238 121519 248240
rect 121453 248235 121519 248238
rect 67725 247752 70226 247754
rect 67725 247696 67730 247752
rect 67786 247696 70226 247752
rect 67725 247694 70226 247696
rect 67725 247691 67791 247694
rect 121637 247618 121703 247621
rect 119876 247616 121703 247618
rect 67633 247210 67699 247213
rect 70166 247210 70226 247588
rect 119876 247560 121642 247616
rect 121698 247560 121703 247616
rect 119876 247558 121703 247560
rect 121637 247555 121703 247558
rect 67633 247208 70226 247210
rect 67633 247152 67638 247208
rect 67694 247152 70226 247208
rect 67633 247150 70226 247152
rect 67633 247147 67699 247150
rect 121545 246938 121611 246941
rect 119876 246936 121611 246938
rect 70166 246394 70226 246908
rect 119876 246880 121550 246936
rect 121606 246880 121611 246936
rect 119876 246878 121611 246880
rect 121545 246875 121611 246878
rect 64830 246334 70226 246394
rect 58934 245652 58940 245716
rect 59004 245714 59010 245716
rect 64830 245714 64890 246334
rect 121453 246258 121519 246261
rect 119876 246256 121519 246258
rect 59004 245654 64890 245714
rect 69105 245714 69171 245717
rect 70166 245714 70226 246228
rect 119876 246200 121458 246256
rect 121514 246200 121519 246256
rect 119876 246198 121519 246200
rect 121453 246195 121519 246198
rect 69105 245712 70226 245714
rect 69105 245656 69110 245712
rect 69166 245656 70226 245712
rect 69105 245654 70226 245656
rect 59004 245652 59010 245654
rect 69105 245651 69171 245654
rect 121637 245578 121703 245581
rect 119876 245576 121703 245578
rect 67633 245306 67699 245309
rect 70350 245306 70410 245548
rect 119876 245520 121642 245576
rect 121698 245520 121703 245576
rect 119876 245518 121703 245520
rect 121637 245515 121703 245518
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 67633 245304 70410 245306
rect 67633 245248 67638 245304
rect 67694 245248 70410 245304
rect 67633 245246 70410 245248
rect 67633 245243 67699 245246
rect 121729 244898 121795 244901
rect 119876 244896 121795 244898
rect 68093 244354 68159 244357
rect 70166 244354 70226 244868
rect 119876 244840 121734 244896
rect 121790 244840 121795 244896
rect 119876 244838 121795 244840
rect 121729 244835 121795 244838
rect 68093 244352 70226 244354
rect 68093 244296 68098 244352
rect 68154 244296 70226 244352
rect 68093 244294 70226 244296
rect 68093 244291 68159 244294
rect 121545 244218 121611 244221
rect 119876 244216 121611 244218
rect 69197 243674 69263 243677
rect 70350 243674 70410 244188
rect 119876 244160 121550 244216
rect 121606 244160 121611 244216
rect 119876 244158 121611 244160
rect 121545 244155 121611 244158
rect 69197 243672 70410 243674
rect 69197 243616 69202 243672
rect 69258 243616 70410 243672
rect 69197 243614 70410 243616
rect 69197 243611 69263 243614
rect 121453 243538 121519 243541
rect 119876 243536 121519 243538
rect 67633 243266 67699 243269
rect 70350 243266 70410 243508
rect 119876 243480 121458 243536
rect 121514 243480 121519 243536
rect 119876 243478 121519 243480
rect 121453 243475 121519 243478
rect 67633 243264 70410 243266
rect 67633 243208 67638 243264
rect 67694 243208 70410 243264
rect 67633 243206 70410 243208
rect 67633 243203 67699 243206
rect 121453 242858 121519 242861
rect 119876 242856 121519 242858
rect 70166 242314 70226 242828
rect 119876 242800 121458 242856
rect 121514 242800 121519 242856
rect 119876 242798 121519 242800
rect 121453 242795 121519 242798
rect 64830 242254 70226 242314
rect 59118 241708 59124 241772
rect 59188 241770 59194 241772
rect 64830 241770 64890 242254
rect 121545 242178 121611 242181
rect 119876 242176 121611 242178
rect 67633 241906 67699 241909
rect 70166 241906 70226 242148
rect 119876 242120 121550 242176
rect 121606 242120 121611 242176
rect 119876 242118 121611 242120
rect 121545 242115 121611 242118
rect 67633 241904 70226 241906
rect 67633 241848 67638 241904
rect 67694 241848 70226 241904
rect 67633 241846 70226 241848
rect 67633 241843 67699 241846
rect 59188 241710 64890 241770
rect 59188 241708 59194 241710
rect -960 241090 480 241180
rect 3049 241090 3115 241093
rect -960 241088 3115 241090
rect -960 241032 3054 241088
rect 3110 241032 3115 241088
rect -960 241030 3115 241032
rect -960 240940 480 241030
rect 3049 241027 3115 241030
rect 70166 240954 70226 241468
rect 119478 241226 119538 241468
rect 122925 241226 122991 241229
rect 119478 241224 122991 241226
rect 119478 241168 122930 241224
rect 122986 241168 122991 241224
rect 119478 241166 122991 241168
rect 64830 240894 70226 240954
rect 57830 240348 57836 240412
rect 57900 240410 57906 240412
rect 64830 240410 64890 240894
rect 119286 240892 119292 240956
rect 119356 240954 119362 240956
rect 119478 240954 119538 241166
rect 122925 241163 122991 241166
rect 119356 240894 119538 240954
rect 119356 240892 119362 240894
rect 121453 240818 121519 240821
rect 119876 240816 121519 240818
rect 57900 240350 64890 240410
rect 57900 240348 57906 240350
rect 69749 240274 69815 240277
rect 70166 240274 70226 240788
rect 119876 240760 121458 240816
rect 121514 240760 121519 240816
rect 119876 240758 121519 240760
rect 121453 240755 121519 240758
rect 69749 240272 70226 240274
rect 69749 240216 69754 240272
rect 69810 240216 70226 240272
rect 69749 240214 70226 240216
rect 69749 240211 69815 240214
rect 121453 240138 121519 240141
rect 119876 240136 121519 240138
rect 119876 240080 121458 240136
rect 121514 240080 121519 240136
rect 119876 240078 121519 240080
rect 121453 240075 121519 240078
rect 118734 239804 118740 239868
rect 118804 239866 118810 239868
rect 118957 239866 119023 239869
rect 118804 239864 119023 239866
rect 118804 239808 118962 239864
rect 119018 239808 119023 239864
rect 118804 239806 119023 239808
rect 118804 239804 118810 239806
rect 118957 239803 119023 239806
rect 61745 239458 61811 239461
rect 82077 239458 82143 239461
rect 61745 239456 82143 239458
rect 61745 239400 61750 239456
rect 61806 239400 82082 239456
rect 82138 239400 82143 239456
rect 61745 239398 82143 239400
rect 61745 239395 61811 239398
rect 82077 239395 82143 239398
rect 50981 238642 51047 238645
rect 98361 238642 98427 238645
rect 50981 238640 98427 238642
rect 50981 238584 50986 238640
rect 51042 238584 98366 238640
rect 98422 238584 98427 238640
rect 50981 238582 98427 238584
rect 50981 238579 51047 238582
rect 98361 238579 98427 238582
rect 113817 238642 113883 238645
rect 125726 238642 125732 238644
rect 113817 238640 125732 238642
rect 113817 238584 113822 238640
rect 113878 238584 125732 238640
rect 113817 238582 125732 238584
rect 113817 238579 113883 238582
rect 125726 238580 125732 238582
rect 125796 238580 125802 238644
rect 55029 238506 55095 238509
rect 91921 238506 91987 238509
rect 55029 238504 91987 238506
rect 55029 238448 55034 238504
rect 55090 238448 91926 238504
rect 91982 238448 91987 238504
rect 55029 238446 91987 238448
rect 55029 238443 55095 238446
rect 91921 238443 91987 238446
rect 117037 238506 117103 238509
rect 124254 238506 124260 238508
rect 117037 238504 124260 238506
rect 117037 238448 117042 238504
rect 117098 238448 124260 238504
rect 117037 238446 124260 238448
rect 117037 238443 117103 238446
rect 124254 238444 124260 238446
rect 124324 238444 124330 238508
rect 61878 237220 61884 237284
rect 61948 237282 61954 237284
rect 86217 237282 86283 237285
rect 61948 237280 86283 237282
rect 61948 237224 86222 237280
rect 86278 237224 86283 237280
rect 61948 237222 86283 237224
rect 61948 237220 61954 237222
rect 86217 237219 86283 237222
rect 61694 232460 61700 232524
rect 61764 232522 61770 232524
rect 583017 232522 583083 232525
rect 61764 232520 583083 232522
rect 61764 232464 583022 232520
rect 583078 232464 583083 232520
rect 61764 232462 583083 232464
rect 61764 232460 61770 232462
rect 583017 232459 583083 232462
rect 580533 232386 580599 232389
rect 583520 232386 584960 232476
rect 580533 232384 584960 232386
rect 580533 232328 580538 232384
rect 580594 232328 584960 232384
rect 580533 232326 584960 232328
rect 580533 232323 580599 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 84377 226946 84443 226949
rect 328494 226946 328500 226948
rect 84377 226944 328500 226946
rect 84377 226888 84382 226944
rect 84438 226888 328500 226944
rect 84377 226886 328500 226888
rect 84377 226883 84443 226886
rect 328494 226884 328500 226886
rect 328564 226884 328570 226948
rect 582833 219058 582899 219061
rect 583520 219058 584960 219148
rect 582833 219056 584960 219058
rect 582833 219000 582838 219056
rect 582894 219000 584960 219056
rect 582833 218998 584960 219000
rect 582833 218995 582899 218998
rect 583520 218908 584960 218998
rect 60365 218650 60431 218653
rect 258390 218650 258396 218652
rect 60365 218648 258396 218650
rect 60365 218592 60370 218648
rect 60426 218592 258396 218648
rect 60365 218590 258396 218592
rect 60365 218587 60431 218590
rect 258390 218588 258396 218590
rect 258460 218588 258466 218652
rect 65926 217228 65932 217292
rect 65996 217290 66002 217292
rect 324589 217290 324655 217293
rect 65996 217288 324655 217290
rect 65996 217232 324594 217288
rect 324650 217232 324655 217288
rect 65996 217230 324655 217232
rect 65996 217228 66002 217230
rect 324589 217227 324655 217230
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 52177 211850 52243 211853
rect 262254 211850 262260 211852
rect 52177 211848 262260 211850
rect 52177 211792 52182 211848
rect 52238 211792 262260 211848
rect 52177 211790 262260 211792
rect 52177 211787 52243 211790
rect 262254 211788 262260 211790
rect 262324 211788 262330 211852
rect 49509 206274 49575 206277
rect 336774 206274 336780 206276
rect 49509 206272 336780 206274
rect 49509 206216 49514 206272
rect 49570 206216 336780 206272
rect 49509 206214 336780 206216
rect 49509 206211 49575 206214
rect 336774 206212 336780 206214
rect 336844 206212 336850 206276
rect 580441 205730 580507 205733
rect 583520 205730 584960 205820
rect 580441 205728 584960 205730
rect 580441 205672 580446 205728
rect 580502 205672 584960 205728
rect 580441 205670 584960 205672
rect 580441 205667 580507 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3601 201922 3667 201925
rect -960 201920 3667 201922
rect -960 201864 3606 201920
rect 3662 201864 3667 201920
rect -960 201862 3667 201864
rect -960 201772 480 201862
rect 3601 201859 3667 201862
rect 1301 200698 1367 200701
rect 118918 200698 118924 200700
rect 1301 200696 118924 200698
rect 1301 200640 1306 200696
rect 1362 200640 118924 200696
rect 1301 200638 118924 200640
rect 1301 200635 1367 200638
rect 118918 200636 118924 200638
rect 118988 200636 118994 200700
rect 218697 192538 218763 192541
rect 339718 192538 339724 192540
rect 218697 192536 339724 192538
rect 218697 192480 218702 192536
rect 218758 192480 339724 192536
rect 218697 192478 339724 192480
rect 218697 192475 218763 192478
rect 339718 192476 339724 192478
rect 339788 192476 339794 192540
rect 583109 192538 583175 192541
rect 583520 192538 584960 192628
rect 583109 192536 584960 192538
rect 583109 192480 583114 192536
rect 583170 192480 584960 192536
rect 583109 192478 584960 192480
rect 583109 192475 583175 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 229737 186962 229803 186965
rect 259678 186962 259684 186964
rect 229737 186960 259684 186962
rect 229737 186904 229742 186960
rect 229798 186904 259684 186960
rect 229737 186902 259684 186904
rect 229737 186899 229803 186902
rect 259678 186900 259684 186902
rect 259748 186900 259754 186964
rect 210509 185602 210575 185605
rect 256734 185602 256740 185604
rect 210509 185600 256740 185602
rect 210509 185544 210514 185600
rect 210570 185544 256740 185600
rect 210509 185542 256740 185544
rect 210509 185539 210575 185542
rect 256734 185540 256740 185542
rect 256804 185540 256810 185604
rect 159357 183018 159423 183021
rect 191189 183018 191255 183021
rect 159357 183016 191255 183018
rect 159357 182960 159362 183016
rect 159418 182960 191194 183016
rect 191250 182960 191255 183016
rect 159357 182958 191255 182960
rect 159357 182955 159423 182958
rect 191189 182955 191255 182958
rect 60641 182882 60707 182885
rect 343817 182882 343883 182885
rect 60641 182880 343883 182882
rect 60641 182824 60646 182880
rect 60702 182824 343822 182880
rect 343878 182824 343883 182880
rect 60641 182822 343883 182824
rect 60641 182819 60707 182822
rect 343817 182819 343883 182822
rect 74533 181386 74599 181389
rect 323025 181386 323091 181389
rect 74533 181384 323091 181386
rect 74533 181328 74538 181384
rect 74594 181328 323030 181384
rect 323086 181328 323091 181384
rect 74533 181326 323091 181328
rect 74533 181323 74599 181326
rect 323025 181323 323091 181326
rect 295977 180162 296043 180165
rect 331438 180162 331444 180164
rect 295977 180160 331444 180162
rect 295977 180104 295982 180160
rect 296038 180104 331444 180160
rect 295977 180102 331444 180104
rect 295977 180099 296043 180102
rect 331438 180100 331444 180102
rect 331508 180100 331514 180164
rect 166349 180026 166415 180029
rect 189717 180026 189783 180029
rect 166349 180024 189783 180026
rect 166349 179968 166354 180024
rect 166410 179968 189722 180024
rect 189778 179968 189783 180024
rect 166349 179966 189783 179968
rect 166349 179963 166415 179966
rect 189717 179963 189783 179966
rect 300209 180026 300275 180029
rect 338246 180026 338252 180028
rect 300209 180024 338252 180026
rect 300209 179968 300214 180024
rect 300270 179968 338252 180024
rect 300209 179966 338252 179968
rect 300209 179963 300275 179966
rect 338246 179964 338252 179966
rect 338316 179964 338322 180028
rect 97257 179482 97323 179485
rect 166206 179482 166212 179484
rect 97257 179480 166212 179482
rect 97257 179424 97262 179480
rect 97318 179424 166212 179480
rect 97257 179422 166212 179424
rect 97257 179419 97323 179422
rect 166206 179420 166212 179422
rect 166276 179420 166282 179484
rect 580257 179210 580323 179213
rect 583520 179210 584960 179300
rect 580257 179208 584960 179210
rect 580257 179152 580262 179208
rect 580318 179152 584960 179208
rect 580257 179150 584960 179152
rect 580257 179147 580323 179150
rect 583520 179060 584960 179150
rect 240777 178802 240843 178805
rect 266486 178802 266492 178804
rect 240777 178800 266492 178802
rect 240777 178744 240782 178800
rect 240838 178744 266492 178800
rect 240777 178742 266492 178744
rect 240777 178739 240843 178742
rect 266486 178740 266492 178742
rect 266556 178740 266562 178804
rect 53649 178666 53715 178669
rect 346669 178666 346735 178669
rect 53649 178664 346735 178666
rect 53649 178608 53654 178664
rect 53710 178608 346674 178664
rect 346730 178608 346735 178664
rect 53649 178606 346735 178608
rect 53649 178603 53715 178606
rect 346669 178603 346735 178606
rect 98310 177652 98316 177716
rect 98380 177714 98386 177716
rect 99281 177714 99347 177717
rect 98380 177712 99347 177714
rect 98380 177656 99286 177712
rect 99342 177656 99347 177712
rect 98380 177654 99347 177656
rect 98380 177652 98386 177654
rect 99281 177651 99347 177654
rect 104566 177652 104572 177716
rect 104636 177714 104642 177716
rect 104801 177714 104867 177717
rect 104636 177712 104867 177714
rect 104636 177656 104806 177712
rect 104862 177656 104867 177712
rect 104636 177654 104867 177656
rect 104636 177652 104642 177654
rect 104801 177651 104867 177654
rect 106958 177652 106964 177716
rect 107028 177714 107034 177716
rect 107561 177714 107627 177717
rect 110689 177716 110755 177717
rect 110638 177714 110644 177716
rect 107028 177712 107627 177714
rect 107028 177656 107566 177712
rect 107622 177656 107627 177712
rect 107028 177654 107627 177656
rect 110598 177654 110644 177714
rect 110708 177712 110755 177716
rect 110750 177656 110755 177712
rect 107028 177652 107034 177654
rect 107561 177651 107627 177654
rect 110638 177652 110644 177654
rect 110708 177652 110755 177656
rect 114318 177652 114324 177716
rect 114388 177714 114394 177716
rect 114461 177714 114527 177717
rect 115841 177716 115907 177717
rect 116945 177716 117011 177717
rect 115790 177714 115796 177716
rect 114388 177712 114527 177714
rect 114388 177656 114466 177712
rect 114522 177656 114527 177712
rect 114388 177654 114527 177656
rect 115750 177654 115796 177714
rect 115860 177712 115907 177716
rect 116894 177714 116900 177716
rect 115902 177656 115907 177712
rect 114388 177652 114394 177654
rect 110689 177651 110755 177652
rect 114461 177651 114527 177654
rect 115790 177652 115796 177654
rect 115860 177652 115907 177656
rect 116854 177654 116900 177714
rect 116964 177712 117011 177716
rect 117006 177656 117011 177712
rect 116894 177652 116900 177654
rect 116964 177652 117011 177656
rect 119470 177652 119476 177716
rect 119540 177714 119546 177716
rect 119981 177714 120047 177717
rect 119540 177712 120047 177714
rect 119540 177656 119986 177712
rect 120042 177656 120047 177712
rect 119540 177654 120047 177656
rect 119540 177652 119546 177654
rect 115841 177651 115907 177652
rect 116945 177651 117011 177652
rect 119981 177651 120047 177654
rect 120758 177652 120764 177716
rect 120828 177714 120834 177716
rect 120901 177714 120967 177717
rect 120828 177712 120967 177714
rect 120828 177656 120906 177712
rect 120962 177656 120967 177712
rect 120828 177654 120967 177656
rect 120828 177652 120834 177654
rect 120901 177651 120967 177654
rect 129406 177652 129412 177716
rect 129476 177714 129482 177716
rect 129641 177714 129707 177717
rect 130745 177716 130811 177717
rect 130694 177714 130700 177716
rect 129476 177712 129707 177714
rect 129476 177656 129646 177712
rect 129702 177656 129707 177712
rect 129476 177654 129707 177656
rect 130654 177654 130700 177714
rect 130764 177712 130811 177716
rect 130806 177656 130811 177712
rect 129476 177652 129482 177654
rect 129641 177651 129707 177654
rect 130694 177652 130700 177654
rect 130764 177652 130811 177656
rect 130745 177651 130811 177652
rect 240869 177578 240935 177581
rect 249190 177578 249196 177580
rect 240869 177576 249196 177578
rect 240869 177520 240874 177576
rect 240930 177520 249196 177576
rect 240869 177518 249196 177520
rect 240869 177515 240935 177518
rect 249190 177516 249196 177518
rect 249260 177516 249266 177580
rect 231117 177442 231183 177445
rect 249374 177442 249380 177444
rect 231117 177440 249380 177442
rect 231117 177384 231122 177440
rect 231178 177384 249380 177440
rect 231117 177382 249380 177384
rect 231117 177379 231183 177382
rect 249374 177380 249380 177382
rect 249444 177380 249450 177444
rect 313917 177442 313983 177445
rect 335118 177442 335124 177444
rect 313917 177440 335124 177442
rect 313917 177384 313922 177440
rect 313978 177384 335124 177440
rect 313917 177382 335124 177384
rect 313917 177379 313983 177382
rect 335118 177380 335124 177382
rect 335188 177380 335194 177444
rect 162117 177306 162183 177309
rect 185577 177306 185643 177309
rect 162117 177304 185643 177306
rect 162117 177248 162122 177304
rect 162178 177248 185582 177304
rect 185638 177248 185643 177304
rect 162117 177246 185643 177248
rect 162117 177243 162183 177246
rect 185577 177243 185643 177246
rect 232497 177306 232563 177309
rect 334198 177306 334204 177308
rect 232497 177304 334204 177306
rect 232497 177248 232502 177304
rect 232558 177248 334204 177304
rect 232497 177246 334204 177248
rect 232497 177243 232563 177246
rect 334198 177244 334204 177246
rect 334268 177244 334274 177308
rect 97022 176972 97028 177036
rect 97092 177034 97098 177036
rect 97257 177034 97323 177037
rect 112161 177036 112227 177037
rect 112110 177034 112116 177036
rect 97092 177032 97323 177034
rect 97092 176976 97262 177032
rect 97318 176976 97323 177032
rect 97092 176974 97323 176976
rect 112070 176974 112116 177034
rect 112180 177032 112227 177036
rect 112222 176976 112227 177032
rect 97092 176972 97098 176974
rect 97257 176971 97323 176974
rect 112110 176972 112116 176974
rect 112180 176972 112227 176976
rect 124438 176972 124444 177036
rect 124508 177034 124514 177036
rect 125409 177034 125475 177037
rect 124508 177032 125475 177034
rect 124508 176976 125414 177032
rect 125470 176976 125475 177032
rect 124508 176974 125475 176976
rect 124508 176972 124514 176974
rect 112161 176971 112227 176972
rect 125409 176971 125475 176974
rect 105670 176836 105676 176900
rect 105740 176898 105746 176900
rect 168230 176898 168236 176900
rect 105740 176838 168236 176898
rect 105740 176836 105746 176838
rect 168230 176836 168236 176838
rect 168300 176836 168306 176900
rect 100661 176762 100727 176765
rect 102041 176764 102107 176765
rect 101990 176762 101996 176764
rect 99422 176760 100727 176762
rect 99422 176704 100666 176760
rect 100722 176704 100727 176760
rect 99422 176702 100727 176704
rect 101950 176702 101996 176762
rect 102060 176760 102107 176764
rect 103329 176762 103395 176765
rect 108113 176764 108179 176765
rect 108062 176762 108068 176764
rect 102102 176704 102107 176760
rect 99422 176492 99482 176702
rect 100661 176699 100727 176702
rect 101990 176700 101996 176702
rect 102060 176700 102107 176704
rect 102041 176699 102107 176700
rect 103286 176760 103395 176762
rect 103286 176704 103334 176760
rect 103390 176704 103395 176760
rect 103286 176699 103395 176704
rect 108022 176702 108068 176762
rect 108132 176760 108179 176764
rect 108174 176704 108179 176760
rect 108062 176700 108068 176702
rect 108132 176700 108179 176704
rect 109534 176700 109540 176764
rect 109604 176762 109610 176764
rect 110045 176762 110111 176765
rect 109604 176760 110111 176762
rect 109604 176704 110050 176760
rect 110106 176704 110111 176760
rect 109604 176702 110111 176704
rect 109604 176700 109610 176702
rect 108113 176699 108179 176700
rect 110045 176699 110111 176702
rect 123150 176700 123156 176764
rect 123220 176762 123226 176764
rect 123293 176762 123359 176765
rect 123220 176760 123359 176762
rect 123220 176704 123298 176760
rect 123354 176704 123359 176760
rect 123220 176702 123359 176704
rect 123220 176700 123226 176702
rect 123293 176699 123359 176702
rect 125726 176700 125732 176764
rect 125796 176762 125802 176764
rect 125869 176762 125935 176765
rect 128261 176762 128327 176765
rect 133137 176764 133203 176765
rect 134425 176764 134491 176765
rect 136081 176764 136147 176765
rect 148225 176764 148291 176765
rect 133086 176762 133092 176764
rect 125796 176760 125935 176762
rect 125796 176704 125874 176760
rect 125930 176704 125935 176760
rect 125796 176702 125935 176704
rect 125796 176700 125802 176702
rect 125869 176699 125935 176702
rect 128126 176760 128327 176762
rect 128126 176704 128266 176760
rect 128322 176704 128327 176760
rect 128126 176702 128327 176704
rect 133046 176702 133092 176762
rect 133156 176760 133203 176764
rect 134374 176762 134380 176764
rect 133198 176704 133203 176760
rect 103286 176492 103346 176699
rect 128126 176492 128186 176702
rect 128261 176699 128327 176702
rect 133086 176700 133092 176702
rect 133156 176700 133203 176704
rect 134334 176702 134380 176762
rect 134444 176760 134491 176764
rect 136030 176762 136036 176764
rect 134486 176704 134491 176760
rect 134374 176700 134380 176702
rect 134444 176700 134491 176704
rect 135990 176702 136036 176762
rect 136100 176760 136147 176764
rect 148174 176762 148180 176764
rect 136142 176704 136147 176760
rect 136030 176700 136036 176702
rect 136100 176700 136147 176704
rect 148134 176702 148180 176762
rect 148244 176760 148291 176764
rect 148286 176704 148291 176760
rect 148174 176700 148180 176702
rect 148244 176700 148291 176704
rect 133137 176699 133203 176700
rect 134425 176699 134491 176700
rect 136081 176699 136147 176700
rect 148225 176699 148291 176700
rect 99414 176428 99420 176492
rect 99484 176428 99490 176492
rect 103278 176428 103284 176492
rect 103348 176428 103354 176492
rect 128118 176428 128124 176492
rect 128188 176428 128194 176492
rect 244917 176354 244983 176357
rect 263726 176354 263732 176356
rect 244917 176352 263732 176354
rect 244917 176296 244922 176352
rect 244978 176296 263732 176352
rect 244917 176294 263732 176296
rect 244917 176291 244983 176294
rect 263726 176292 263732 176294
rect 263796 176292 263802 176356
rect 213913 176218 213979 176221
rect 242249 176218 242315 176221
rect 213913 176216 217242 176218
rect 213913 176160 213918 176216
rect 213974 176160 217242 176216
rect 213913 176158 217242 176160
rect 213913 176155 213979 176158
rect -960 175796 480 176036
rect 217182 175644 217242 176158
rect 242249 176216 248338 176218
rect 242249 176160 242254 176216
rect 242310 176160 248338 176216
rect 242249 176158 248338 176160
rect 242249 176155 242315 176158
rect 248278 175644 248338 176158
rect 320817 175946 320883 175949
rect 326061 175946 326127 175949
rect 320817 175944 326127 175946
rect 320817 175888 320822 175944
rect 320878 175888 326066 175944
rect 326122 175888 326127 175944
rect 320817 175886 326127 175888
rect 320817 175883 320883 175886
rect 326061 175883 326127 175886
rect 296069 175810 296135 175813
rect 296069 175808 321386 175810
rect 296069 175752 296074 175808
rect 296130 175752 321386 175808
rect 296069 175750 321386 175752
rect 296069 175747 296135 175750
rect 296670 175614 310132 175674
rect 127065 175540 127131 175541
rect 132033 175540 132099 175541
rect 158897 175540 158963 175541
rect 113214 175476 113220 175540
rect 113284 175538 113290 175540
rect 127014 175538 127020 175540
rect 113284 175478 122850 175538
rect 126974 175478 127020 175538
rect 127084 175536 127131 175540
rect 131982 175538 131988 175540
rect 127126 175480 127131 175536
rect 113284 175476 113290 175478
rect 100753 175404 100819 175405
rect 118417 175404 118483 175405
rect 121913 175404 121979 175405
rect 100702 175402 100708 175404
rect 100662 175342 100708 175402
rect 100772 175400 100819 175404
rect 118366 175402 118372 175404
rect 100814 175344 100819 175400
rect 100702 175340 100708 175342
rect 100772 175340 100819 175344
rect 118326 175342 118372 175402
rect 118436 175400 118483 175404
rect 121862 175402 121868 175404
rect 118478 175344 118483 175400
rect 118366 175340 118372 175342
rect 118436 175340 118483 175344
rect 121822 175342 121868 175402
rect 121932 175400 121979 175404
rect 121974 175344 121979 175400
rect 121862 175340 121868 175342
rect 121932 175340 121979 175344
rect 122790 175402 122850 175478
rect 127014 175476 127020 175478
rect 127084 175476 127131 175480
rect 131942 175478 131988 175538
rect 132052 175536 132099 175540
rect 158846 175538 158852 175540
rect 132094 175480 132099 175536
rect 131982 175476 131988 175478
rect 132052 175476 132099 175480
rect 158806 175478 158852 175538
rect 158916 175536 158963 175540
rect 158958 175480 158963 175536
rect 158846 175476 158852 175478
rect 158916 175476 158963 175480
rect 127065 175475 127131 175476
rect 132033 175475 132099 175476
rect 158897 175475 158963 175476
rect 166390 175402 166396 175404
rect 122790 175342 166396 175402
rect 166390 175340 166396 175342
rect 166460 175340 166466 175404
rect 262070 175340 262076 175404
rect 262140 175402 262146 175404
rect 296670 175402 296730 175614
rect 321326 175508 321386 175750
rect 262140 175342 296730 175402
rect 262140 175340 262146 175342
rect 100753 175339 100819 175340
rect 118417 175339 118483 175340
rect 121913 175339 121979 175340
rect 249241 175266 249307 175269
rect 248952 175264 249307 175266
rect 248952 175208 249246 175264
rect 249302 175208 249307 175264
rect 248952 175206 249307 175208
rect 249241 175203 249307 175206
rect 306966 175204 306972 175268
rect 307036 175266 307042 175268
rect 321461 175266 321527 175269
rect 307036 175206 310040 175266
rect 321461 175264 321570 175266
rect 321461 175208 321466 175264
rect 321522 175208 321570 175264
rect 307036 175204 307042 175206
rect 321461 175203 321570 175208
rect 213913 175130 213979 175133
rect 213913 175128 217242 175130
rect 213913 175072 213918 175128
rect 213974 175072 217242 175128
rect 213913 175070 217242 175072
rect 213913 175067 213979 175070
rect 217182 174964 217242 175070
rect 307477 174858 307543 174861
rect 307477 174856 310040 174858
rect 307477 174800 307482 174856
rect 307538 174800 310040 174856
rect 307477 174798 310040 174800
rect 307477 174795 307543 174798
rect 214005 174722 214071 174725
rect 249190 174722 249196 174724
rect 214005 174720 217242 174722
rect 214005 174664 214010 174720
rect 214066 174664 217242 174720
rect 214005 174662 217242 174664
rect 248952 174662 249196 174722
rect 214005 174659 214071 174662
rect 217182 174284 217242 174662
rect 249190 174660 249196 174662
rect 249260 174660 249266 174724
rect 321510 174692 321570 175203
rect 307569 174450 307635 174453
rect 307569 174448 310040 174450
rect 307569 174392 307574 174448
rect 307630 174392 310040 174448
rect 307569 174390 310040 174392
rect 307569 174387 307635 174390
rect 249149 174314 249215 174317
rect 248952 174312 249215 174314
rect 248952 174256 249154 174312
rect 249210 174256 249215 174312
rect 248952 174254 249215 174256
rect 249149 174251 249215 174254
rect 307661 174042 307727 174045
rect 324313 174042 324379 174045
rect 307661 174040 310040 174042
rect 307661 173984 307666 174040
rect 307722 173984 310040 174040
rect 307661 173982 310040 173984
rect 321908 174040 324379 174042
rect 321908 173984 324318 174040
rect 324374 173984 324379 174040
rect 321908 173982 324379 173984
rect 307661 173979 307727 173982
rect 324313 173979 324379 173982
rect 213913 173770 213979 173773
rect 252461 173770 252527 173773
rect 213913 173768 217242 173770
rect 213913 173712 213918 173768
rect 213974 173712 217242 173768
rect 213913 173710 217242 173712
rect 248952 173768 252527 173770
rect 248952 173712 252466 173768
rect 252522 173712 252527 173768
rect 248952 173710 252527 173712
rect 213913 173707 213979 173710
rect 217182 173604 217242 173710
rect 252461 173707 252527 173710
rect 307569 173634 307635 173637
rect 307569 173632 310040 173634
rect 307569 173576 307574 173632
rect 307630 173576 310040 173632
rect 307569 173574 310040 173576
rect 307569 173571 307635 173574
rect 214649 173362 214715 173365
rect 249374 173362 249380 173364
rect 214649 173360 217242 173362
rect 214649 173304 214654 173360
rect 214710 173304 217242 173360
rect 214649 173302 217242 173304
rect 248952 173302 249380 173362
rect 214649 173299 214715 173302
rect 217182 172924 217242 173302
rect 249374 173300 249380 173302
rect 249444 173300 249450 173364
rect 307477 173226 307543 173229
rect 324313 173226 324379 173229
rect 307477 173224 310040 173226
rect 307477 173168 307482 173224
rect 307538 173168 310040 173224
rect 307477 173166 310040 173168
rect 321908 173224 324379 173226
rect 321908 173168 324318 173224
rect 324374 173168 324379 173224
rect 321908 173166 324379 173168
rect 307477 173163 307543 173166
rect 324313 173163 324379 173166
rect 249149 172818 249215 172821
rect 248952 172816 249215 172818
rect 248952 172760 249154 172816
rect 249210 172760 249215 172816
rect 248952 172758 249215 172760
rect 249149 172755 249215 172758
rect 307661 172682 307727 172685
rect 307661 172680 310040 172682
rect 307661 172624 307666 172680
rect 307722 172624 310040 172680
rect 307661 172622 310040 172624
rect 307661 172619 307727 172622
rect 213913 172410 213979 172413
rect 249333 172410 249399 172413
rect 324405 172410 324471 172413
rect 213913 172408 217242 172410
rect 213913 172352 213918 172408
rect 213974 172352 217242 172408
rect 213913 172350 217242 172352
rect 248952 172408 249399 172410
rect 248952 172352 249338 172408
rect 249394 172352 249399 172408
rect 248952 172350 249399 172352
rect 321908 172408 324471 172410
rect 321908 172352 324410 172408
rect 324466 172352 324471 172408
rect 321908 172350 324471 172352
rect 213913 172347 213979 172350
rect 217182 172244 217242 172350
rect 249333 172347 249399 172350
rect 324405 172347 324471 172350
rect 306557 172274 306623 172277
rect 306557 172272 310040 172274
rect 306557 172216 306562 172272
rect 306618 172216 310040 172272
rect 306557 172214 310040 172216
rect 306557 172211 306623 172214
rect 214005 172002 214071 172005
rect 214005 172000 217242 172002
rect 214005 171944 214010 172000
rect 214066 171944 217242 172000
rect 214005 171942 217242 171944
rect 214005 171939 214071 171942
rect 167821 171594 167887 171597
rect 164694 171592 167887 171594
rect 164694 171536 167826 171592
rect 167882 171536 167887 171592
rect 217182 171564 217242 171942
rect 252645 171866 252711 171869
rect 248952 171864 252711 171866
rect 248952 171808 252650 171864
rect 252706 171808 252711 171864
rect 248952 171806 252711 171808
rect 252645 171803 252711 171806
rect 307569 171866 307635 171869
rect 307569 171864 310040 171866
rect 307569 171808 307574 171864
rect 307630 171808 310040 171864
rect 307569 171806 310040 171808
rect 307569 171803 307635 171806
rect 164694 171534 167887 171536
rect 167821 171531 167887 171534
rect 252461 171458 252527 171461
rect 248952 171456 252527 171458
rect 248952 171400 252466 171456
rect 252522 171400 252527 171456
rect 248952 171398 252527 171400
rect 252461 171395 252527 171398
rect 307661 171458 307727 171461
rect 307661 171456 310040 171458
rect 307661 171400 307666 171456
rect 307722 171400 310040 171456
rect 307661 171398 310040 171400
rect 307661 171395 307727 171398
rect 321878 171186 321938 171700
rect 326061 171186 326127 171189
rect 216998 171126 217242 171186
rect 321878 171184 326127 171186
rect 321878 171128 326066 171184
rect 326122 171128 326127 171184
rect 321878 171126 326127 171128
rect 216998 171050 217058 171126
rect 215250 170990 217058 171050
rect 217182 171020 217242 171126
rect 326061 171123 326127 171126
rect 307293 171050 307359 171053
rect 307293 171048 310040 171050
rect 307293 170992 307298 171048
rect 307354 170992 310040 171048
rect 307293 170990 310040 170992
rect 214465 170914 214531 170917
rect 215250 170914 215310 170990
rect 307293 170987 307359 170990
rect 252461 170914 252527 170917
rect 324313 170914 324379 170917
rect 214465 170912 215310 170914
rect 214465 170856 214470 170912
rect 214526 170856 215310 170912
rect 214465 170854 215310 170856
rect 248952 170912 252527 170914
rect 248952 170856 252466 170912
rect 252522 170856 252527 170912
rect 248952 170854 252527 170856
rect 321908 170912 324379 170914
rect 321908 170856 324318 170912
rect 324374 170856 324379 170912
rect 321908 170854 324379 170856
rect 214465 170851 214531 170854
rect 252461 170851 252527 170854
rect 324313 170851 324379 170854
rect 214925 170778 214991 170781
rect 214925 170776 217242 170778
rect 214925 170720 214930 170776
rect 214986 170720 217242 170776
rect 214925 170718 217242 170720
rect 214925 170715 214991 170718
rect 217182 170340 217242 170718
rect 307661 170642 307727 170645
rect 307661 170640 310040 170642
rect 307661 170584 307666 170640
rect 307722 170584 310040 170640
rect 307661 170582 310040 170584
rect 307661 170579 307727 170582
rect 252277 170506 252343 170509
rect 248952 170504 252343 170506
rect 248952 170448 252282 170504
rect 252338 170448 252343 170504
rect 248952 170446 252343 170448
rect 252277 170443 252343 170446
rect 307477 170234 307543 170237
rect 307477 170232 310040 170234
rect 307477 170176 307482 170232
rect 307538 170176 310040 170232
rect 307477 170174 310040 170176
rect 307477 170171 307543 170174
rect 252369 170098 252435 170101
rect 323209 170098 323275 170101
rect 248952 170096 252435 170098
rect 248952 170040 252374 170096
rect 252430 170040 252435 170096
rect 248952 170038 252435 170040
rect 321908 170096 323275 170098
rect 321908 170040 323214 170096
rect 323270 170040 323275 170096
rect 321908 170038 323275 170040
rect 252369 170035 252435 170038
rect 323209 170035 323275 170038
rect 307385 169826 307451 169829
rect 216998 169766 217242 169826
rect 213913 169690 213979 169693
rect 216998 169690 217058 169766
rect 213913 169688 217058 169690
rect 213913 169632 213918 169688
rect 213974 169632 217058 169688
rect 217182 169660 217242 169766
rect 307385 169824 310040 169826
rect 307385 169768 307390 169824
rect 307446 169768 310040 169824
rect 307385 169766 310040 169768
rect 307385 169763 307451 169766
rect 321277 169690 321343 169693
rect 321277 169688 321386 169690
rect 213913 169630 217058 169632
rect 321277 169632 321282 169688
rect 321338 169632 321386 169688
rect 213913 169627 213979 169630
rect 321277 169627 321386 169632
rect 252461 169554 252527 169557
rect 248952 169552 252527 169554
rect 248952 169496 252466 169552
rect 252522 169496 252527 169552
rect 248952 169494 252527 169496
rect 252461 169491 252527 169494
rect 214005 169418 214071 169421
rect 214005 169416 217242 169418
rect 214005 169360 214010 169416
rect 214066 169360 217242 169416
rect 321326 169388 321386 169627
rect 214005 169358 217242 169360
rect 214005 169355 214071 169358
rect 217182 168980 217242 169358
rect 307569 169282 307635 169285
rect 307569 169280 310040 169282
rect 307569 169224 307574 169280
rect 307630 169224 310040 169280
rect 307569 169222 310040 169224
rect 307569 169219 307635 169222
rect 252369 169146 252435 169149
rect 248952 169144 252435 169146
rect 248952 169088 252374 169144
rect 252430 169088 252435 169144
rect 248952 169086 252435 169088
rect 252369 169083 252435 169086
rect 307661 168874 307727 168877
rect 307661 168872 310040 168874
rect 307661 168816 307666 168872
rect 307722 168816 310040 168872
rect 307661 168814 310040 168816
rect 307661 168811 307727 168814
rect 252461 168602 252527 168605
rect 324313 168602 324379 168605
rect 248952 168600 252527 168602
rect 248952 168544 252466 168600
rect 252522 168544 252527 168600
rect 248952 168542 252527 168544
rect 321908 168600 324379 168602
rect 321908 168544 324318 168600
rect 324374 168544 324379 168600
rect 321908 168542 324379 168544
rect 252461 168539 252527 168542
rect 324313 168539 324379 168542
rect 307109 168466 307175 168469
rect 216998 168406 217242 168466
rect 213913 168330 213979 168333
rect 216998 168330 217058 168406
rect 213913 168328 217058 168330
rect 213913 168272 213918 168328
rect 213974 168272 217058 168328
rect 217182 168300 217242 168406
rect 307109 168464 310040 168466
rect 307109 168408 307114 168464
rect 307170 168408 310040 168464
rect 307109 168406 310040 168408
rect 307109 168403 307175 168406
rect 213913 168270 217058 168272
rect 213913 168267 213979 168270
rect 252461 168194 252527 168197
rect 248952 168192 252527 168194
rect 248952 168136 252466 168192
rect 252522 168136 252527 168192
rect 248952 168134 252527 168136
rect 252461 168131 252527 168134
rect 214005 168058 214071 168061
rect 307293 168058 307359 168061
rect 214005 168056 217242 168058
rect 214005 168000 214010 168056
rect 214066 168000 217242 168056
rect 214005 167998 217242 168000
rect 214005 167995 214071 167998
rect 217182 167620 217242 167998
rect 307293 168056 310040 168058
rect 307293 168000 307298 168056
rect 307354 168000 310040 168056
rect 307293 167998 310040 168000
rect 307293 167995 307359 167998
rect 324313 167786 324379 167789
rect 321908 167784 324379 167786
rect 321908 167728 324318 167784
rect 324374 167728 324379 167784
rect 321908 167726 324379 167728
rect 324313 167723 324379 167726
rect 252461 167650 252527 167653
rect 248952 167648 252527 167650
rect 248952 167592 252466 167648
rect 252522 167592 252527 167648
rect 248952 167590 252527 167592
rect 252461 167587 252527 167590
rect 307477 167650 307543 167653
rect 307477 167648 310040 167650
rect 307477 167592 307482 167648
rect 307538 167592 310040 167648
rect 307477 167590 310040 167592
rect 307477 167587 307543 167590
rect 252369 167242 252435 167245
rect 248952 167240 252435 167242
rect 248952 167184 252374 167240
rect 252430 167184 252435 167240
rect 248952 167182 252435 167184
rect 252369 167179 252435 167182
rect 307661 167242 307727 167245
rect 307661 167240 310040 167242
rect 307661 167184 307666 167240
rect 307722 167184 310040 167240
rect 307661 167182 310040 167184
rect 307661 167179 307727 167182
rect 324405 167106 324471 167109
rect 321908 167104 324471 167106
rect 321908 167048 324410 167104
rect 324466 167048 324471 167104
rect 321908 167046 324471 167048
rect 324405 167043 324471 167046
rect 214741 166970 214807 166973
rect 216998 166970 217242 167010
rect 214741 166968 217242 166970
rect 214741 166912 214746 166968
rect 214802 166950 217242 166968
rect 214802 166912 217058 166950
rect 217182 166940 217242 166950
rect 214741 166910 217058 166912
rect 214741 166907 214807 166910
rect 307569 166834 307635 166837
rect 307569 166832 310040 166834
rect 307569 166776 307574 166832
rect 307630 166776 310040 166832
rect 307569 166774 310040 166776
rect 307569 166771 307635 166774
rect 214005 166698 214071 166701
rect 249793 166698 249859 166701
rect 214005 166696 217242 166698
rect 214005 166640 214010 166696
rect 214066 166640 217242 166696
rect 214005 166638 217242 166640
rect 248952 166696 249859 166698
rect 248952 166640 249798 166696
rect 249854 166640 249859 166696
rect 248952 166638 249859 166640
rect 214005 166635 214071 166638
rect 217182 166396 217242 166638
rect 249793 166635 249859 166638
rect 307109 166426 307175 166429
rect 307109 166424 310040 166426
rect 307109 166368 307114 166424
rect 307170 166368 310040 166424
rect 307109 166366 310040 166368
rect 307109 166363 307175 166366
rect 252461 166290 252527 166293
rect 324313 166290 324379 166293
rect 248952 166288 252527 166290
rect 248952 166232 252466 166288
rect 252522 166232 252527 166288
rect 248952 166230 252527 166232
rect 321908 166288 324379 166290
rect 321908 166232 324318 166288
rect 324374 166232 324379 166288
rect 321908 166230 324379 166232
rect 252461 166227 252527 166230
rect 324313 166227 324379 166230
rect 213913 166154 213979 166157
rect 213913 166152 217242 166154
rect 213913 166096 213918 166152
rect 213974 166096 217242 166152
rect 213913 166094 217242 166096
rect 213913 166091 213979 166094
rect 217182 165716 217242 166094
rect 307661 165882 307727 165885
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 307661 165880 310040 165882
rect 307661 165824 307666 165880
rect 307722 165824 310040 165880
rect 307661 165822 310040 165824
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 307661 165819 307727 165822
rect 580165 165819 580231 165822
rect 252369 165746 252435 165749
rect 248952 165744 252435 165746
rect 248952 165688 252374 165744
rect 252430 165688 252435 165744
rect 583520 165732 584960 165822
rect 248952 165686 252435 165688
rect 252369 165683 252435 165686
rect 307017 165474 307083 165477
rect 324313 165474 324379 165477
rect 307017 165472 310040 165474
rect 307017 165416 307022 165472
rect 307078 165416 310040 165472
rect 307017 165414 310040 165416
rect 321908 165472 324379 165474
rect 321908 165416 324318 165472
rect 324374 165416 324379 165472
rect 321908 165414 324379 165416
rect 307017 165411 307083 165414
rect 324313 165411 324379 165414
rect 213913 165338 213979 165341
rect 252461 165338 252527 165341
rect 213913 165336 217242 165338
rect 213913 165280 213918 165336
rect 213974 165280 217242 165336
rect 213913 165278 217242 165280
rect 248952 165336 252527 165338
rect 248952 165280 252466 165336
rect 252522 165280 252527 165336
rect 248952 165278 252527 165280
rect 213913 165275 213979 165278
rect 217182 165036 217242 165278
rect 252461 165275 252527 165278
rect 307109 165066 307175 165069
rect 307109 165064 310040 165066
rect 307109 165008 307114 165064
rect 307170 165008 310040 165064
rect 307109 165006 310040 165008
rect 307109 165003 307175 165006
rect 214005 164794 214071 164797
rect 252369 164794 252435 164797
rect 324405 164794 324471 164797
rect 214005 164792 217242 164794
rect 214005 164736 214010 164792
rect 214066 164736 217242 164792
rect 214005 164734 217242 164736
rect 248952 164792 252435 164794
rect 248952 164736 252374 164792
rect 252430 164736 252435 164792
rect 248952 164734 252435 164736
rect 321908 164792 324471 164794
rect 321908 164736 324410 164792
rect 324466 164736 324471 164792
rect 321908 164734 324471 164736
rect 214005 164731 214071 164734
rect 217182 164356 217242 164734
rect 252369 164731 252435 164734
rect 324405 164731 324471 164734
rect 307201 164658 307267 164661
rect 307201 164656 310040 164658
rect 307201 164600 307206 164656
rect 307262 164600 310040 164656
rect 307201 164598 310040 164600
rect 307201 164595 307267 164598
rect 251357 164386 251423 164389
rect 248952 164384 251423 164386
rect 248952 164328 251362 164384
rect 251418 164328 251423 164384
rect 248952 164326 251423 164328
rect 251357 164323 251423 164326
rect 307661 164250 307727 164253
rect 307661 164248 310040 164250
rect 307661 164192 307666 164248
rect 307722 164192 310040 164248
rect 307661 164190 310040 164192
rect 307661 164187 307727 164190
rect 252369 163978 252435 163981
rect 324313 163978 324379 163981
rect 248952 163976 252435 163978
rect 248952 163920 252374 163976
rect 252430 163920 252435 163976
rect 248952 163918 252435 163920
rect 321908 163976 324379 163978
rect 321908 163920 324318 163976
rect 324374 163920 324379 163976
rect 321908 163918 324379 163920
rect 252369 163915 252435 163918
rect 324313 163915 324379 163918
rect 307569 163842 307635 163845
rect 200070 163782 217242 163842
rect 166390 163100 166396 163164
rect 166460 163162 166466 163164
rect 200070 163162 200130 163782
rect 217182 163676 217242 163782
rect 307569 163840 310040 163842
rect 307569 163784 307574 163840
rect 307630 163784 310040 163840
rect 307569 163782 310040 163784
rect 307569 163779 307635 163782
rect 213913 163434 213979 163437
rect 252461 163434 252527 163437
rect 213913 163432 217426 163434
rect 213913 163376 213918 163432
rect 213974 163376 217426 163432
rect 213913 163374 217426 163376
rect 248952 163432 252527 163434
rect 248952 163376 252466 163432
rect 252522 163376 252527 163432
rect 248952 163374 252527 163376
rect 213913 163371 213979 163374
rect 166460 163102 200130 163162
rect 166460 163100 166466 163102
rect 217366 162996 217426 163374
rect 252461 163371 252527 163374
rect 306741 163434 306807 163437
rect 306741 163432 310040 163434
rect 306741 163376 306746 163432
rect 306802 163376 310040 163432
rect 306741 163374 310040 163376
rect 306741 163371 306807 163374
rect 324405 163162 324471 163165
rect 321908 163160 324471 163162
rect 321908 163104 324410 163160
rect 324466 163104 324471 163160
rect 321908 163102 324471 163104
rect 324405 163099 324471 163102
rect 252277 163026 252343 163029
rect 248952 163024 252343 163026
rect -960 162890 480 162980
rect 248952 162968 252282 163024
rect 252338 162968 252343 163024
rect 248952 162966 252343 162968
rect 252277 162963 252343 162966
rect 307661 163026 307727 163029
rect 307661 163024 310040 163026
rect 307661 162968 307666 163024
rect 307722 162968 310040 163024
rect 307661 162966 310040 162968
rect 307661 162963 307727 162966
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 213913 162618 213979 162621
rect 213913 162616 217242 162618
rect 213913 162560 213918 162616
rect 213974 162560 217242 162616
rect 213913 162558 217242 162560
rect 213913 162555 213979 162558
rect 217182 162316 217242 162558
rect 252553 162482 252619 162485
rect 248952 162480 252619 162482
rect 248952 162424 252558 162480
rect 252614 162424 252619 162480
rect 248952 162422 252619 162424
rect 252553 162419 252619 162422
rect 307477 162482 307543 162485
rect 324313 162482 324379 162485
rect 307477 162480 310040 162482
rect 307477 162424 307482 162480
rect 307538 162424 310040 162480
rect 307477 162422 310040 162424
rect 321908 162480 324379 162482
rect 321908 162424 324318 162480
rect 324374 162424 324379 162480
rect 321908 162422 324379 162424
rect 307477 162419 307543 162422
rect 324313 162419 324379 162422
rect 214005 162074 214071 162077
rect 307569 162074 307635 162077
rect 214005 162072 217242 162074
rect 214005 162016 214010 162072
rect 214066 162016 217242 162072
rect 307569 162072 310040 162074
rect 214005 162014 217242 162016
rect 214005 162011 214071 162014
rect 217182 161772 217242 162014
rect 248860 161970 249442 162030
rect 307569 162016 307574 162072
rect 307630 162016 310040 162072
rect 307569 162014 310040 162016
rect 307569 162011 307635 162014
rect 249382 161802 249442 161970
rect 262254 161802 262260 161804
rect 249382 161742 262260 161802
rect 262254 161740 262260 161742
rect 262324 161740 262330 161804
rect 307661 161666 307727 161669
rect 324405 161666 324471 161669
rect 307661 161664 310040 161666
rect 307661 161608 307666 161664
rect 307722 161608 310040 161664
rect 307661 161606 310040 161608
rect 321908 161664 324471 161666
rect 321908 161608 324410 161664
rect 324466 161608 324471 161664
rect 321908 161606 324471 161608
rect 307661 161603 307727 161606
rect 324405 161603 324471 161606
rect 252461 161530 252527 161533
rect 248952 161528 252527 161530
rect 248952 161472 252466 161528
rect 252522 161472 252527 161528
rect 248952 161470 252527 161472
rect 252461 161467 252527 161470
rect 214649 161258 214715 161261
rect 306557 161258 306623 161261
rect 214649 161256 217242 161258
rect 214649 161200 214654 161256
rect 214710 161200 217242 161256
rect 214649 161198 217242 161200
rect 214649 161195 214715 161198
rect 217182 161092 217242 161198
rect 306557 161256 310040 161258
rect 306557 161200 306562 161256
rect 306618 161200 310040 161256
rect 306557 161198 310040 161200
rect 306557 161195 306623 161198
rect 252461 161122 252527 161125
rect 248952 161120 252527 161122
rect 248952 161064 252466 161120
rect 252522 161064 252527 161120
rect 248952 161062 252527 161064
rect 252461 161059 252527 161062
rect 213913 160850 213979 160853
rect 307661 160850 307727 160853
rect 324313 160850 324379 160853
rect 213913 160848 217242 160850
rect 213913 160792 213918 160848
rect 213974 160792 217242 160848
rect 213913 160790 217242 160792
rect 213913 160787 213979 160790
rect 217182 160412 217242 160790
rect 307661 160848 310040 160850
rect 307661 160792 307666 160848
rect 307722 160792 310040 160848
rect 307661 160790 310040 160792
rect 321908 160848 324379 160850
rect 321908 160792 324318 160848
rect 324374 160792 324379 160848
rect 321908 160790 324379 160792
rect 307661 160787 307727 160790
rect 324313 160787 324379 160790
rect 252369 160578 252435 160581
rect 248952 160576 252435 160578
rect 248952 160520 252374 160576
rect 252430 160520 252435 160576
rect 248952 160518 252435 160520
rect 252369 160515 252435 160518
rect 307569 160442 307635 160445
rect 307569 160440 310040 160442
rect 307569 160384 307574 160440
rect 307630 160384 310040 160440
rect 307569 160382 310040 160384
rect 307569 160379 307635 160382
rect 252001 160170 252067 160173
rect 324405 160170 324471 160173
rect 248952 160168 252067 160170
rect 248952 160112 252006 160168
rect 252062 160112 252067 160168
rect 248952 160110 252067 160112
rect 321908 160168 324471 160170
rect 321908 160112 324410 160168
rect 324466 160112 324471 160168
rect 321908 160110 324471 160112
rect 252001 160107 252067 160110
rect 324405 160107 324471 160110
rect 307569 160034 307635 160037
rect 307569 160032 310040 160034
rect 307569 159976 307574 160032
rect 307630 159976 310040 160032
rect 307569 159974 310040 159976
rect 307569 159971 307635 159974
rect 321737 159898 321803 159901
rect 321694 159896 321803 159898
rect 321694 159840 321742 159896
rect 321798 159840 321803 159896
rect 321694 159835 321803 159840
rect 217182 159218 217242 159732
rect 251265 159626 251331 159629
rect 248952 159624 251331 159626
rect 248952 159568 251270 159624
rect 251326 159568 251331 159624
rect 248952 159566 251331 159568
rect 251265 159563 251331 159566
rect 307109 159626 307175 159629
rect 307109 159624 310040 159626
rect 307109 159568 307114 159624
rect 307170 159568 310040 159624
rect 307109 159566 310040 159568
rect 307109 159563 307175 159566
rect 250621 159354 250687 159357
rect 258390 159354 258396 159356
rect 250621 159352 258396 159354
rect 250621 159296 250626 159352
rect 250682 159296 258396 159352
rect 250621 159294 258396 159296
rect 250621 159291 250687 159294
rect 258390 159292 258396 159294
rect 258460 159292 258466 159356
rect 321694 159324 321754 159835
rect 252461 159218 252527 159221
rect 200070 159158 217242 159218
rect 248952 159216 252527 159218
rect 248952 159160 252466 159216
rect 252522 159160 252527 159216
rect 248952 159158 252527 159160
rect 168230 158748 168236 158812
rect 168300 158810 168306 158812
rect 200070 158810 200130 159158
rect 252461 159155 252527 159158
rect 307661 159082 307727 159085
rect 307661 159080 310040 159082
rect 168300 158750 200130 158810
rect 213913 158810 213979 158813
rect 217366 158810 217426 159052
rect 307661 159024 307666 159080
rect 307722 159024 310040 159080
rect 307661 159022 310040 159024
rect 307661 159019 307727 159022
rect 251449 158810 251515 158813
rect 213913 158808 217426 158810
rect 213913 158752 213918 158808
rect 213974 158752 217426 158808
rect 213913 158750 217426 158752
rect 248952 158808 251515 158810
rect 248952 158752 251454 158808
rect 251510 158752 251515 158808
rect 248952 158750 251515 158752
rect 168300 158748 168306 158750
rect 213913 158747 213979 158750
rect 251449 158747 251515 158750
rect 213913 158674 213979 158677
rect 252001 158674 252067 158677
rect 259678 158674 259684 158676
rect 213913 158672 217242 158674
rect 213913 158616 213918 158672
rect 213974 158616 217242 158672
rect 213913 158614 217242 158616
rect 213913 158611 213979 158614
rect 217182 158372 217242 158614
rect 252001 158672 259684 158674
rect 252001 158616 252006 158672
rect 252062 158616 259684 158672
rect 252001 158614 259684 158616
rect 252001 158611 252067 158614
rect 259678 158612 259684 158614
rect 259748 158612 259754 158676
rect 306925 158674 306991 158677
rect 306925 158672 310040 158674
rect 306925 158616 306930 158672
rect 306986 158616 310040 158672
rect 306925 158614 310040 158616
rect 306925 158611 306991 158614
rect 324313 158538 324379 158541
rect 321908 158536 324379 158538
rect 321908 158480 324318 158536
rect 324374 158480 324379 158536
rect 321908 158478 324379 158480
rect 324313 158475 324379 158478
rect 252461 158266 252527 158269
rect 248952 158264 252527 158266
rect 248952 158208 252466 158264
rect 252522 158208 252527 158264
rect 248952 158206 252527 158208
rect 252461 158203 252527 158206
rect 307569 158266 307635 158269
rect 307569 158264 310040 158266
rect 307569 158208 307574 158264
rect 307630 158208 310040 158264
rect 307569 158206 310040 158208
rect 307569 158203 307635 158206
rect 214005 158130 214071 158133
rect 214005 158128 217242 158130
rect 214005 158072 214010 158128
rect 214066 158072 217242 158128
rect 214005 158070 217242 158072
rect 214005 158067 214071 158070
rect 217182 157692 217242 158070
rect 251173 157858 251239 157861
rect 248952 157856 251239 157858
rect 248952 157800 251178 157856
rect 251234 157800 251239 157856
rect 248952 157798 251239 157800
rect 251173 157795 251239 157798
rect 307661 157858 307727 157861
rect 324405 157858 324471 157861
rect 307661 157856 310040 157858
rect 307661 157800 307666 157856
rect 307722 157800 310040 157856
rect 307661 157798 310040 157800
rect 321908 157856 324471 157858
rect 321908 157800 324410 157856
rect 324466 157800 324471 157856
rect 321908 157798 324471 157800
rect 307661 157795 307727 157798
rect 324405 157795 324471 157798
rect 307385 157450 307451 157453
rect 307385 157448 310040 157450
rect 307385 157392 307390 157448
rect 307446 157392 310040 157448
rect 307385 157390 310040 157392
rect 307385 157387 307451 157390
rect 213913 157314 213979 157317
rect 213913 157312 217242 157314
rect 213913 157256 213918 157312
rect 213974 157256 217242 157312
rect 213913 157254 217242 157256
rect 213913 157251 213979 157254
rect 217182 157148 217242 157254
rect 248860 157210 249442 157270
rect 249382 157178 249442 157210
rect 263726 157178 263732 157180
rect 249382 157118 263732 157178
rect 263726 157116 263732 157118
rect 263796 157116 263802 157180
rect 307477 157042 307543 157045
rect 324313 157042 324379 157045
rect 307477 157040 310040 157042
rect 307477 156984 307482 157040
rect 307538 156984 310040 157040
rect 307477 156982 310040 156984
rect 321908 157040 324379 157042
rect 321908 156984 324318 157040
rect 324374 156984 324379 157040
rect 321908 156982 324379 156984
rect 307477 156979 307543 156982
rect 324313 156979 324379 156982
rect 214005 156906 214071 156909
rect 252461 156906 252527 156909
rect 214005 156904 217242 156906
rect 214005 156848 214010 156904
rect 214066 156848 217242 156904
rect 214005 156846 217242 156848
rect 248952 156904 252527 156906
rect 248952 156848 252466 156904
rect 252522 156848 252527 156904
rect 248952 156846 252527 156848
rect 214005 156843 214071 156846
rect 217182 156468 217242 156846
rect 252461 156843 252527 156846
rect 307569 156634 307635 156637
rect 307569 156632 310040 156634
rect 307569 156576 307574 156632
rect 307630 156576 310040 156632
rect 307569 156574 310040 156576
rect 307569 156571 307635 156574
rect 252369 156362 252435 156365
rect 324313 156362 324379 156365
rect 248952 156360 252435 156362
rect 248952 156304 252374 156360
rect 252430 156304 252435 156360
rect 248952 156302 252435 156304
rect 321908 156360 324379 156362
rect 321908 156304 324318 156360
rect 324374 156304 324379 156360
rect 321908 156302 324379 156304
rect 252369 156299 252435 156302
rect 324313 156299 324379 156302
rect 307661 156226 307727 156229
rect 307661 156224 310040 156226
rect 307661 156168 307666 156224
rect 307722 156168 310040 156224
rect 307661 156166 310040 156168
rect 307661 156163 307727 156166
rect 213913 155954 213979 155957
rect 252461 155954 252527 155957
rect 213913 155952 217242 155954
rect 213913 155896 213918 155952
rect 213974 155896 217242 155952
rect 213913 155894 217242 155896
rect 248952 155952 252527 155954
rect 248952 155896 252466 155952
rect 252522 155896 252527 155952
rect 248952 155894 252527 155896
rect 213913 155891 213979 155894
rect 217182 155788 217242 155894
rect 252461 155891 252527 155894
rect 306557 155682 306623 155685
rect 306557 155680 310040 155682
rect 306557 155624 306562 155680
rect 306618 155624 310040 155680
rect 306557 155622 310040 155624
rect 306557 155619 306623 155622
rect 324313 155546 324379 155549
rect 321908 155544 324379 155546
rect 321908 155488 324318 155544
rect 324374 155488 324379 155544
rect 321908 155486 324379 155488
rect 324313 155483 324379 155486
rect 251541 155410 251607 155413
rect 248952 155408 251607 155410
rect 248952 155352 251546 155408
rect 251602 155352 251607 155408
rect 248952 155350 251607 155352
rect 251541 155347 251607 155350
rect 307661 155274 307727 155277
rect 307661 155272 310040 155274
rect 307661 155216 307666 155272
rect 307722 155216 310040 155272
rect 307661 155214 310040 155216
rect 307661 155211 307727 155214
rect 166206 154532 166212 154596
rect 166276 154594 166282 154596
rect 217182 154594 217242 155108
rect 252461 155002 252527 155005
rect 248952 155000 252527 155002
rect 248952 154944 252466 155000
rect 252522 154944 252527 155000
rect 248952 154942 252527 154944
rect 252461 154939 252527 154942
rect 307201 154866 307267 154869
rect 307201 154864 310040 154866
rect 307201 154808 307206 154864
rect 307262 154808 310040 154864
rect 307201 154806 310040 154808
rect 307201 154803 307267 154806
rect 324405 154730 324471 154733
rect 321908 154728 324471 154730
rect 321908 154672 324410 154728
rect 324466 154672 324471 154728
rect 321908 154670 324471 154672
rect 324405 154667 324471 154670
rect 166276 154534 217242 154594
rect 166276 154532 166282 154534
rect 252829 154458 252895 154461
rect 248952 154456 252895 154458
rect 214005 153914 214071 153917
rect 217182 153914 217242 154428
rect 248952 154400 252834 154456
rect 252890 154400 252895 154456
rect 248952 154398 252895 154400
rect 252829 154395 252895 154398
rect 306557 154458 306623 154461
rect 306557 154456 310040 154458
rect 306557 154400 306562 154456
rect 306618 154400 310040 154456
rect 306557 154398 310040 154400
rect 306557 154395 306623 154398
rect 252461 154050 252527 154053
rect 248952 154048 252527 154050
rect 248952 153992 252466 154048
rect 252522 153992 252527 154048
rect 248952 153990 252527 153992
rect 252461 153987 252527 153990
rect 307569 154050 307635 154053
rect 324313 154050 324379 154053
rect 307569 154048 310040 154050
rect 307569 153992 307574 154048
rect 307630 153992 310040 154048
rect 307569 153990 310040 153992
rect 321908 154048 324379 154050
rect 321908 153992 324318 154048
rect 324374 153992 324379 154048
rect 321908 153990 324379 153992
rect 307569 153987 307635 153990
rect 324313 153987 324379 153990
rect 214005 153912 217242 153914
rect 214005 153856 214010 153912
rect 214066 153856 217242 153912
rect 214005 153854 217242 153856
rect 214005 153851 214071 153854
rect 213913 153506 213979 153509
rect 217182 153506 217242 153748
rect 307661 153642 307727 153645
rect 307661 153640 310040 153642
rect 307661 153584 307666 153640
rect 307722 153584 310040 153640
rect 307661 153582 310040 153584
rect 307661 153579 307727 153582
rect 249885 153506 249951 153509
rect 213913 153504 217242 153506
rect 213913 153448 213918 153504
rect 213974 153448 217242 153504
rect 213913 153446 217242 153448
rect 248952 153504 249951 153506
rect 248952 153448 249890 153504
rect 249946 153448 249951 153504
rect 248952 153446 249951 153448
rect 213913 153443 213979 153446
rect 249885 153443 249951 153446
rect 306649 153234 306715 153237
rect 324313 153234 324379 153237
rect 306649 153232 310040 153234
rect 306649 153176 306654 153232
rect 306710 153176 310040 153232
rect 306649 153174 310040 153176
rect 321908 153232 324379 153234
rect 321908 153176 324318 153232
rect 324374 153176 324379 153232
rect 321908 153174 324379 153176
rect 306649 153171 306715 153174
rect 324313 153171 324379 153174
rect 252461 153098 252527 153101
rect 248952 153096 252527 153098
rect 214005 152690 214071 152693
rect 217182 152690 217242 153068
rect 248952 153040 252466 153096
rect 252522 153040 252527 153096
rect 248952 153038 252527 153040
rect 252461 153035 252527 153038
rect 252369 152690 252435 152693
rect 214005 152688 217242 152690
rect 214005 152632 214010 152688
rect 214066 152632 217242 152688
rect 214005 152630 217242 152632
rect 248952 152688 252435 152690
rect 248952 152632 252374 152688
rect 252430 152632 252435 152688
rect 248952 152630 252435 152632
rect 214005 152627 214071 152630
rect 252369 152627 252435 152630
rect 306557 152690 306623 152693
rect 580349 152690 580415 152693
rect 583520 152690 584960 152780
rect 306557 152688 310040 152690
rect 306557 152632 306562 152688
rect 306618 152632 310040 152688
rect 306557 152630 310040 152632
rect 580349 152688 584960 152690
rect 580349 152632 580354 152688
rect 580410 152632 584960 152688
rect 580349 152630 584960 152632
rect 306557 152627 306623 152630
rect 580349 152627 580415 152630
rect 583520 152540 584960 152630
rect 213913 152010 213979 152013
rect 217182 152010 217242 152524
rect 324405 152418 324471 152421
rect 321908 152416 324471 152418
rect 321908 152360 324410 152416
rect 324466 152360 324471 152416
rect 321908 152358 324471 152360
rect 324405 152355 324471 152358
rect 307477 152282 307543 152285
rect 307477 152280 310040 152282
rect 307477 152224 307482 152280
rect 307538 152224 310040 152280
rect 307477 152222 310040 152224
rect 307477 152219 307543 152222
rect 255262 152146 255268 152148
rect 248952 152086 255268 152146
rect 255262 152084 255268 152086
rect 255332 152084 255338 152148
rect 213913 152008 217242 152010
rect 213913 151952 213918 152008
rect 213974 151952 217242 152008
rect 213913 151950 217242 151952
rect 213913 151947 213979 151950
rect 214557 151874 214623 151877
rect 307661 151874 307727 151877
rect 214557 151872 217058 151874
rect 214557 151816 214562 151872
rect 214618 151830 217058 151872
rect 307661 151872 310040 151874
rect 217182 151830 217242 151844
rect 214618 151816 217242 151830
rect 214557 151814 217242 151816
rect 214557 151811 214623 151814
rect 216998 151770 217242 151814
rect 307661 151816 307666 151872
rect 307722 151816 310040 151872
rect 307661 151814 310040 151816
rect 307661 151811 307727 151814
rect 252369 151738 252435 151741
rect 324313 151738 324379 151741
rect 248952 151736 252435 151738
rect 248952 151680 252374 151736
rect 252430 151680 252435 151736
rect 248952 151678 252435 151680
rect 321908 151736 324379 151738
rect 321908 151680 324318 151736
rect 324374 151680 324379 151736
rect 321908 151678 324379 151680
rect 252369 151675 252435 151678
rect 324313 151675 324379 151678
rect 307477 151466 307543 151469
rect 307477 151464 310040 151466
rect 307477 151408 307482 151464
rect 307538 151408 310040 151464
rect 307477 151406 310040 151408
rect 307477 151403 307543 151406
rect 252461 151194 252527 151197
rect 248952 151192 252527 151194
rect 214741 150786 214807 150789
rect 217182 150786 217242 151164
rect 248952 151136 252466 151192
rect 252522 151136 252527 151192
rect 248952 151134 252527 151136
rect 252461 151131 252527 151134
rect 307661 151058 307727 151061
rect 307661 151056 310040 151058
rect 307661 151000 307666 151056
rect 307722 151000 310040 151056
rect 307661 150998 310040 151000
rect 307661 150995 307727 150998
rect 323117 150922 323183 150925
rect 321908 150920 323183 150922
rect 321908 150864 323122 150920
rect 323178 150864 323183 150920
rect 321908 150862 323183 150864
rect 323117 150859 323183 150862
rect 251357 150786 251423 150789
rect 214741 150784 217242 150786
rect 214741 150728 214746 150784
rect 214802 150728 217242 150784
rect 214741 150726 217242 150728
rect 248952 150784 251423 150786
rect 248952 150728 251362 150784
rect 251418 150728 251423 150784
rect 248952 150726 251423 150728
rect 214741 150723 214807 150726
rect 251357 150723 251423 150726
rect 213913 150650 213979 150653
rect 307569 150650 307635 150653
rect 213913 150648 217242 150650
rect 213913 150592 213918 150648
rect 213974 150592 217242 150648
rect 213913 150590 217242 150592
rect 213913 150587 213979 150590
rect 217182 150484 217242 150590
rect 307569 150648 310040 150650
rect 307569 150592 307574 150648
rect 307630 150592 310040 150648
rect 307569 150590 310040 150592
rect 307569 150587 307635 150590
rect 252461 150242 252527 150245
rect 248952 150240 252527 150242
rect 248952 150184 252466 150240
rect 252522 150184 252527 150240
rect 248952 150182 252527 150184
rect 252461 150179 252527 150182
rect 307477 150242 307543 150245
rect 307477 150240 310040 150242
rect 307477 150184 307482 150240
rect 307538 150184 310040 150240
rect 307477 150182 310040 150184
rect 307477 150179 307543 150182
rect 214005 150106 214071 150109
rect 324313 150106 324379 150109
rect 214005 150104 217242 150106
rect 214005 150048 214010 150104
rect 214066 150048 217242 150104
rect 214005 150046 217242 150048
rect 321908 150104 324379 150106
rect 321908 150048 324318 150104
rect 324374 150048 324379 150104
rect 321908 150046 324379 150048
rect 214005 150043 214071 150046
rect -960 149834 480 149924
rect 3509 149834 3575 149837
rect -960 149832 3575 149834
rect -960 149776 3514 149832
rect 3570 149776 3575 149832
rect 217182 149804 217242 150046
rect 324313 150043 324379 150046
rect 252093 149834 252159 149837
rect 248952 149832 252159 149834
rect -960 149774 3575 149776
rect 248952 149776 252098 149832
rect 252154 149776 252159 149832
rect 248952 149774 252159 149776
rect -960 149684 480 149774
rect 3509 149771 3575 149774
rect 252093 149771 252159 149774
rect 306557 149834 306623 149837
rect 306557 149832 310040 149834
rect 306557 149776 306562 149832
rect 306618 149776 310040 149832
rect 306557 149774 310040 149776
rect 306557 149771 306623 149774
rect 214649 149562 214715 149565
rect 214649 149560 217242 149562
rect 214649 149504 214654 149560
rect 214710 149504 217242 149560
rect 214649 149502 217242 149504
rect 214649 149499 214715 149502
rect 217182 149124 217242 149502
rect 324405 149426 324471 149429
rect 321908 149424 324471 149426
rect 321908 149368 324410 149424
rect 324466 149368 324471 149424
rect 321908 149366 324471 149368
rect 324405 149363 324471 149366
rect 252277 149290 252343 149293
rect 248952 149288 252343 149290
rect 248952 149232 252282 149288
rect 252338 149232 252343 149288
rect 248952 149230 252343 149232
rect 252277 149227 252343 149230
rect 307569 149290 307635 149293
rect 307569 149288 310040 149290
rect 307569 149232 307574 149288
rect 307630 149232 310040 149288
rect 307569 149230 310040 149232
rect 307569 149227 307635 149230
rect 252461 148882 252527 148885
rect 248952 148880 252527 148882
rect 248952 148824 252466 148880
rect 252522 148824 252527 148880
rect 248952 148822 252527 148824
rect 252461 148819 252527 148822
rect 307293 148882 307359 148885
rect 307293 148880 310040 148882
rect 307293 148824 307298 148880
rect 307354 148824 310040 148880
rect 307293 148822 310040 148824
rect 307293 148819 307359 148822
rect 213913 148746 213979 148749
rect 213913 148744 217242 148746
rect 213913 148688 213918 148744
rect 213974 148688 217242 148744
rect 213913 148686 217242 148688
rect 213913 148683 213979 148686
rect 217182 148444 217242 148686
rect 324313 148610 324379 148613
rect 321908 148608 324379 148610
rect 321908 148552 324318 148608
rect 324374 148552 324379 148608
rect 321908 148550 324379 148552
rect 324313 148547 324379 148550
rect 307661 148474 307727 148477
rect 307661 148472 310040 148474
rect 307661 148416 307666 148472
rect 307722 148416 310040 148472
rect 307661 148414 310040 148416
rect 307661 148411 307727 148414
rect 252369 148338 252435 148341
rect 248952 148336 252435 148338
rect 248952 148280 252374 148336
rect 252430 148280 252435 148336
rect 248952 148278 252435 148280
rect 252369 148275 252435 148278
rect 213913 148066 213979 148069
rect 213913 148064 217242 148066
rect 213913 148008 213918 148064
rect 213974 148008 217242 148064
rect 213913 148006 217242 148008
rect 213913 148003 213979 148006
rect 217182 147900 217242 148006
rect 309550 147962 310132 148022
rect 252277 147930 252343 147933
rect 248952 147928 252343 147930
rect 248952 147872 252282 147928
rect 252338 147872 252343 147928
rect 248952 147870 252343 147872
rect 252277 147867 252343 147870
rect 305637 147794 305703 147797
rect 309550 147794 309610 147962
rect 325877 147794 325943 147797
rect 305637 147792 309610 147794
rect 305637 147736 305642 147792
rect 305698 147736 309610 147792
rect 305637 147734 309610 147736
rect 321908 147792 325943 147794
rect 321908 147736 325882 147792
rect 325938 147736 325943 147792
rect 321908 147734 325943 147736
rect 305637 147731 305703 147734
rect 325877 147731 325943 147734
rect 307385 147658 307451 147661
rect 307385 147656 310040 147658
rect 307385 147600 307390 147656
rect 307446 147600 310040 147656
rect 307385 147598 310040 147600
rect 307385 147595 307451 147598
rect 256734 147522 256740 147524
rect 248952 147462 256740 147522
rect 256734 147460 256740 147462
rect 256804 147460 256810 147524
rect 307293 147250 307359 147253
rect 307293 147248 310040 147250
rect 214005 146706 214071 146709
rect 217182 146706 217242 147220
rect 307293 147192 307298 147248
rect 307354 147192 310040 147248
rect 307293 147190 310040 147192
rect 307293 147187 307359 147190
rect 324313 147114 324379 147117
rect 321908 147112 324379 147114
rect 321908 147056 324318 147112
rect 324374 147056 324379 147112
rect 321908 147054 324379 147056
rect 324313 147051 324379 147054
rect 252737 146978 252803 146981
rect 248952 146976 252803 146978
rect 248952 146920 252742 146976
rect 252798 146920 252803 146976
rect 248952 146918 252803 146920
rect 252737 146915 252803 146918
rect 306925 146842 306991 146845
rect 306925 146840 310040 146842
rect 306925 146784 306930 146840
rect 306986 146784 310040 146840
rect 306925 146782 310040 146784
rect 306925 146779 306991 146782
rect 214005 146704 217242 146706
rect 214005 146648 214010 146704
rect 214066 146648 217242 146704
rect 214005 146646 217242 146648
rect 214005 146643 214071 146646
rect 252461 146570 252527 146573
rect 248952 146568 252527 146570
rect 213913 146434 213979 146437
rect 213913 146432 216874 146434
rect 213913 146376 213918 146432
rect 213974 146376 216874 146432
rect 213913 146374 216874 146376
rect 213913 146371 213979 146374
rect 216814 146298 216874 146374
rect 217366 146298 217426 146540
rect 248952 146512 252466 146568
rect 252522 146512 252527 146568
rect 248952 146510 252527 146512
rect 252461 146507 252527 146510
rect 306741 146434 306807 146437
rect 306741 146432 310040 146434
rect 306741 146376 306746 146432
rect 306802 146376 310040 146432
rect 306741 146374 310040 146376
rect 306741 146371 306807 146374
rect 324313 146298 324379 146301
rect 216814 146238 217426 146298
rect 321908 146296 324379 146298
rect 321908 146240 324318 146296
rect 324374 146240 324379 146296
rect 321908 146238 324379 146240
rect 324313 146235 324379 146238
rect 252461 146026 252527 146029
rect 248952 146024 252527 146026
rect 248952 145968 252466 146024
rect 252522 145968 252527 146024
rect 248952 145966 252527 145968
rect 252461 145963 252527 145966
rect 307569 145890 307635 145893
rect 307569 145888 310040 145890
rect 214005 145346 214071 145349
rect 217182 145346 217242 145860
rect 307569 145832 307574 145888
rect 307630 145832 310040 145888
rect 307569 145830 310040 145832
rect 307569 145827 307635 145830
rect 252369 145618 252435 145621
rect 248952 145616 252435 145618
rect 248952 145560 252374 145616
rect 252430 145560 252435 145616
rect 248952 145558 252435 145560
rect 252369 145555 252435 145558
rect 307477 145482 307543 145485
rect 324313 145482 324379 145485
rect 307477 145480 310040 145482
rect 307477 145424 307482 145480
rect 307538 145424 310040 145480
rect 307477 145422 310040 145424
rect 321908 145480 324379 145482
rect 321908 145424 324318 145480
rect 324374 145424 324379 145480
rect 321908 145422 324379 145424
rect 307477 145419 307543 145422
rect 324313 145419 324379 145422
rect 214005 145344 217242 145346
rect 214005 145288 214010 145344
rect 214066 145288 217242 145344
rect 214005 145286 217242 145288
rect 214005 145283 214071 145286
rect 213913 144938 213979 144941
rect 217366 144938 217426 145180
rect 252277 145074 252343 145077
rect 248952 145072 252343 145074
rect 248952 145016 252282 145072
rect 252338 145016 252343 145072
rect 248952 145014 252343 145016
rect 252277 145011 252343 145014
rect 307661 145074 307727 145077
rect 307661 145072 310040 145074
rect 307661 145016 307666 145072
rect 307722 145016 310040 145072
rect 307661 145014 310040 145016
rect 307661 145011 307727 145014
rect 213913 144936 217426 144938
rect 213913 144880 213918 144936
rect 213974 144880 217426 144936
rect 213913 144878 217426 144880
rect 213913 144875 213979 144878
rect 324313 144802 324379 144805
rect 321908 144800 324379 144802
rect 321908 144744 324318 144800
rect 324374 144744 324379 144800
rect 321908 144742 324379 144744
rect 324313 144739 324379 144742
rect 252185 144666 252251 144669
rect 248952 144664 252251 144666
rect 248952 144608 252190 144664
rect 252246 144608 252251 144664
rect 248952 144606 252251 144608
rect 252185 144603 252251 144606
rect 306557 144666 306623 144669
rect 306557 144664 310040 144666
rect 306557 144608 306562 144664
rect 306618 144608 310040 144664
rect 306557 144606 310040 144608
rect 306557 144603 306623 144606
rect 213913 143986 213979 143989
rect 217182 143986 217242 144500
rect 307661 144258 307727 144261
rect 307661 144256 310040 144258
rect 307661 144200 307666 144256
rect 307722 144200 310040 144256
rect 307661 144198 310040 144200
rect 307661 144195 307727 144198
rect 252461 144122 252527 144125
rect 248952 144120 252527 144122
rect 248952 144064 252466 144120
rect 252522 144064 252527 144120
rect 248952 144062 252527 144064
rect 252461 144059 252527 144062
rect 324405 143986 324471 143989
rect 213913 143984 217242 143986
rect 213913 143928 213918 143984
rect 213974 143928 217242 143984
rect 213913 143926 217242 143928
rect 321908 143984 324471 143986
rect 321908 143928 324410 143984
rect 324466 143928 324471 143984
rect 321908 143926 324471 143928
rect 213913 143923 213979 143926
rect 324405 143923 324471 143926
rect 306649 143850 306715 143853
rect 306649 143848 310040 143850
rect 214833 143578 214899 143581
rect 217182 143578 217242 143820
rect 306649 143792 306654 143848
rect 306710 143792 310040 143848
rect 306649 143790 310040 143792
rect 306649 143787 306715 143790
rect 252369 143714 252435 143717
rect 248952 143712 252435 143714
rect 248952 143656 252374 143712
rect 252430 143656 252435 143712
rect 248952 143654 252435 143656
rect 252369 143651 252435 143654
rect 214833 143576 217242 143578
rect 214833 143520 214838 143576
rect 214894 143520 217242 143576
rect 214833 143518 217242 143520
rect 214833 143515 214899 143518
rect 307569 143442 307635 143445
rect 307569 143440 310040 143442
rect 307569 143384 307574 143440
rect 307630 143384 310040 143440
rect 307569 143382 310040 143384
rect 307569 143379 307635 143382
rect 214005 142762 214071 142765
rect 217182 142762 217242 143276
rect 252461 143170 252527 143173
rect 324313 143170 324379 143173
rect 248952 143168 252527 143170
rect 248952 143112 252466 143168
rect 252522 143112 252527 143168
rect 248952 143110 252527 143112
rect 321908 143168 324379 143170
rect 321908 143112 324318 143168
rect 324374 143112 324379 143168
rect 321908 143110 324379 143112
rect 252461 143107 252527 143110
rect 324313 143107 324379 143110
rect 307661 143034 307727 143037
rect 307661 143032 310040 143034
rect 307661 142976 307666 143032
rect 307722 142976 310040 143032
rect 307661 142974 310040 142976
rect 307661 142971 307727 142974
rect 251633 142762 251699 142765
rect 214005 142760 217242 142762
rect 214005 142704 214010 142760
rect 214066 142704 217242 142760
rect 214005 142702 217242 142704
rect 248952 142760 251699 142762
rect 248952 142704 251638 142760
rect 251694 142704 251699 142760
rect 248952 142702 251699 142704
rect 214005 142699 214071 142702
rect 251633 142699 251699 142702
rect 251766 142700 251772 142764
rect 251836 142762 251842 142764
rect 306741 142762 306807 142765
rect 251836 142760 306807 142762
rect 251836 142704 306746 142760
rect 306802 142704 306807 142760
rect 251836 142702 306807 142704
rect 251836 142700 251842 142702
rect 306741 142699 306807 142702
rect 213913 142354 213979 142357
rect 217182 142354 217242 142596
rect 306465 142490 306531 142493
rect 324405 142490 324471 142493
rect 306465 142488 310040 142490
rect 306465 142432 306470 142488
rect 306526 142432 310040 142488
rect 306465 142430 310040 142432
rect 321908 142488 324471 142490
rect 321908 142432 324410 142488
rect 324466 142432 324471 142488
rect 321908 142430 324471 142432
rect 306465 142427 306531 142430
rect 324405 142427 324471 142430
rect 213913 142352 217242 142354
rect 213913 142296 213918 142352
rect 213974 142296 217242 142352
rect 213913 142294 217242 142296
rect 213913 142291 213979 142294
rect 252369 142218 252435 142221
rect 248952 142216 252435 142218
rect 248952 142160 252374 142216
rect 252430 142160 252435 142216
rect 248952 142158 252435 142160
rect 252369 142155 252435 142158
rect 307201 142082 307267 142085
rect 307201 142080 310040 142082
rect 307201 142024 307206 142080
rect 307262 142024 310040 142080
rect 307201 142022 310040 142024
rect 307201 142019 307267 142022
rect 213913 141402 213979 141405
rect 217182 141402 217242 141916
rect 248860 141706 249442 141766
rect 249382 141538 249442 141706
rect 253197 141674 253263 141677
rect 307109 141674 307175 141677
rect 324313 141674 324379 141677
rect 253197 141672 253674 141674
rect 253197 141616 253202 141672
rect 253258 141616 253674 141672
rect 253197 141614 253674 141616
rect 253197 141611 253263 141614
rect 249382 141478 253490 141538
rect 252461 141402 252527 141405
rect 213913 141400 217242 141402
rect 213913 141344 213918 141400
rect 213974 141344 217242 141400
rect 213913 141342 217242 141344
rect 248952 141400 252527 141402
rect 248952 141344 252466 141400
rect 252522 141344 252527 141400
rect 248952 141342 252527 141344
rect 213913 141339 213979 141342
rect 252461 141339 252527 141342
rect 214005 140994 214071 140997
rect 217182 140994 217242 141236
rect 253430 141130 253490 141478
rect 253614 141402 253674 141614
rect 307109 141672 310040 141674
rect 307109 141616 307114 141672
rect 307170 141616 310040 141672
rect 307109 141614 310040 141616
rect 321908 141672 324379 141674
rect 321908 141616 324318 141672
rect 324374 141616 324379 141672
rect 321908 141614 324379 141616
rect 307109 141611 307175 141614
rect 324313 141611 324379 141614
rect 254526 141476 254532 141540
rect 254596 141538 254602 141540
rect 306649 141538 306715 141541
rect 254596 141536 306715 141538
rect 254596 141480 306654 141536
rect 306710 141480 306715 141536
rect 254596 141478 306715 141480
rect 254596 141476 254602 141478
rect 306649 141475 306715 141478
rect 306966 141402 306972 141404
rect 253614 141342 306972 141402
rect 306966 141340 306972 141342
rect 307036 141340 307042 141404
rect 307518 141204 307524 141268
rect 307588 141266 307594 141268
rect 307588 141206 310040 141266
rect 307588 141204 307594 141206
rect 266486 141130 266492 141132
rect 253430 141070 266492 141130
rect 266486 141068 266492 141070
rect 266556 141068 266562 141132
rect 214005 140992 217242 140994
rect 214005 140936 214010 140992
rect 214066 140936 217242 140992
rect 214005 140934 217242 140936
rect 214005 140931 214071 140934
rect 252369 140858 252435 140861
rect 248952 140856 252435 140858
rect 248952 140800 252374 140856
rect 252430 140800 252435 140856
rect 248952 140798 252435 140800
rect 252369 140795 252435 140798
rect 307385 140858 307451 140861
rect 324497 140858 324563 140861
rect 307385 140856 310040 140858
rect 307385 140800 307390 140856
rect 307446 140800 310040 140856
rect 307385 140798 310040 140800
rect 321908 140856 324563 140858
rect 321908 140800 324502 140856
rect 324558 140800 324563 140856
rect 321908 140798 324563 140800
rect 307385 140795 307451 140798
rect 324497 140795 324563 140798
rect 213269 140042 213335 140045
rect 217182 140042 217242 140556
rect 252001 140450 252067 140453
rect 248952 140448 252067 140450
rect 248952 140392 252006 140448
rect 252062 140392 252067 140448
rect 248952 140390 252067 140392
rect 252001 140387 252067 140390
rect 307661 140450 307727 140453
rect 307661 140448 310040 140450
rect 307661 140392 307666 140448
rect 307722 140392 310040 140448
rect 307661 140390 310040 140392
rect 307661 140387 307727 140390
rect 324313 140178 324379 140181
rect 321908 140176 324379 140178
rect 321908 140120 324318 140176
rect 324374 140120 324379 140176
rect 321908 140118 324379 140120
rect 324313 140115 324379 140118
rect 213269 140040 217242 140042
rect 213269 139984 213274 140040
rect 213330 139984 217242 140040
rect 213269 139982 217242 139984
rect 213269 139979 213335 139982
rect 309504 139938 310132 139998
rect 252461 139906 252527 139909
rect 248952 139904 252527 139906
rect 213913 139498 213979 139501
rect 217182 139498 217242 139876
rect 248952 139848 252466 139904
rect 252522 139848 252527 139904
rect 248952 139846 252527 139848
rect 252461 139843 252527 139846
rect 302734 139708 302740 139772
rect 302804 139770 302810 139772
rect 309504 139770 309564 139938
rect 302804 139710 309564 139770
rect 302804 139708 302810 139710
rect 307293 139634 307359 139637
rect 307293 139632 310040 139634
rect 307293 139576 307298 139632
rect 307354 139576 310040 139632
rect 307293 139574 310040 139576
rect 307293 139571 307359 139574
rect 252369 139498 252435 139501
rect 213913 139496 217242 139498
rect 213913 139440 213918 139496
rect 213974 139440 217242 139496
rect 213913 139438 217242 139440
rect 248952 139496 252435 139498
rect 248952 139440 252374 139496
rect 252430 139440 252435 139496
rect 248952 139438 252435 139440
rect 213913 139435 213979 139438
rect 252369 139435 252435 139438
rect 324313 139362 324379 139365
rect 321908 139360 324379 139362
rect 321908 139304 324318 139360
rect 324374 139304 324379 139360
rect 321908 139302 324379 139304
rect 324313 139299 324379 139302
rect 580206 139300 580212 139364
rect 580276 139362 580282 139364
rect 583520 139362 584960 139452
rect 580276 139302 584960 139362
rect 580276 139300 580282 139302
rect 583520 139212 584960 139302
rect 217182 138818 217242 139196
rect 307569 139090 307635 139093
rect 307569 139088 310040 139090
rect 307569 139032 307574 139088
rect 307630 139032 310040 139088
rect 307569 139030 310040 139032
rect 307569 139027 307635 139030
rect 252461 138954 252527 138957
rect 248952 138952 252527 138954
rect 248952 138896 252466 138952
rect 252522 138896 252527 138952
rect 248952 138894 252527 138896
rect 252461 138891 252527 138894
rect 200070 138758 217242 138818
rect 170438 138076 170444 138140
rect 170508 138138 170514 138140
rect 200070 138138 200130 138758
rect 307661 138682 307727 138685
rect 307661 138680 310040 138682
rect 170508 138078 200130 138138
rect 213913 138138 213979 138141
rect 217182 138138 217242 138652
rect 307661 138624 307666 138680
rect 307722 138624 310040 138680
rect 307661 138622 310040 138624
rect 307661 138619 307727 138622
rect 252369 138546 252435 138549
rect 324497 138546 324563 138549
rect 248952 138544 252435 138546
rect 248952 138488 252374 138544
rect 252430 138488 252435 138544
rect 248952 138486 252435 138488
rect 321908 138544 324563 138546
rect 321908 138488 324502 138544
rect 324558 138488 324563 138544
rect 321908 138486 324563 138488
rect 252369 138483 252435 138486
rect 324497 138483 324563 138486
rect 307293 138274 307359 138277
rect 307293 138272 310040 138274
rect 307293 138216 307298 138272
rect 307354 138216 310040 138272
rect 307293 138214 310040 138216
rect 307293 138211 307359 138214
rect 213913 138136 217242 138138
rect 213913 138080 213918 138136
rect 213974 138080 217242 138136
rect 213913 138078 217242 138080
rect 170508 138076 170514 138078
rect 213913 138075 213979 138078
rect 252502 138002 252508 138004
rect 214465 137458 214531 137461
rect 217182 137458 217242 137972
rect 248952 137942 252508 138002
rect 252502 137940 252508 137942
rect 252572 137940 252578 138004
rect 307569 137866 307635 137869
rect 324313 137866 324379 137869
rect 307569 137864 310040 137866
rect 307569 137808 307574 137864
rect 307630 137808 310040 137864
rect 307569 137806 310040 137808
rect 321908 137864 324379 137866
rect 321908 137808 324318 137864
rect 324374 137808 324379 137864
rect 321908 137806 324379 137808
rect 307569 137803 307635 137806
rect 324313 137803 324379 137806
rect 252461 137594 252527 137597
rect 248952 137592 252527 137594
rect 248952 137536 252466 137592
rect 252522 137536 252527 137592
rect 248952 137534 252527 137536
rect 252461 137531 252527 137534
rect 214465 137456 217242 137458
rect 214465 137400 214470 137456
rect 214526 137400 217242 137456
rect 214465 137398 217242 137400
rect 307661 137458 307727 137461
rect 307661 137456 310040 137458
rect 307661 137400 307666 137456
rect 307722 137400 310040 137456
rect 307661 137398 310040 137400
rect 214465 137395 214531 137398
rect 307661 137395 307727 137398
rect -960 136778 480 136868
rect 2773 136778 2839 136781
rect -960 136776 2839 136778
rect -960 136720 2778 136776
rect 2834 136720 2839 136776
rect -960 136718 2839 136720
rect -960 136628 480 136718
rect 2773 136715 2839 136718
rect 213913 136778 213979 136781
rect 217182 136778 217242 137292
rect 252369 137050 252435 137053
rect 248952 137048 252435 137050
rect 248952 136992 252374 137048
rect 252430 136992 252435 137048
rect 248952 136990 252435 136992
rect 252369 136987 252435 136990
rect 307201 137050 307267 137053
rect 324497 137050 324563 137053
rect 307201 137048 310040 137050
rect 307201 136992 307206 137048
rect 307262 136992 310040 137048
rect 307201 136990 310040 136992
rect 321908 137048 324563 137050
rect 321908 136992 324502 137048
rect 324558 136992 324563 137048
rect 321908 136990 324563 136992
rect 307201 136987 307267 136990
rect 324497 136987 324563 136990
rect 213913 136776 217242 136778
rect 213913 136720 213918 136776
rect 213974 136720 217242 136776
rect 213913 136718 217242 136720
rect 213913 136715 213979 136718
rect 250621 136642 250687 136645
rect 248952 136640 250687 136642
rect 214741 136098 214807 136101
rect 217182 136098 217242 136612
rect 248952 136584 250626 136640
rect 250682 136584 250687 136640
rect 248952 136582 250687 136584
rect 250621 136579 250687 136582
rect 307477 136642 307543 136645
rect 307477 136640 310040 136642
rect 307477 136584 307482 136640
rect 307538 136584 310040 136640
rect 307477 136582 310040 136584
rect 307477 136579 307543 136582
rect 324313 136370 324379 136373
rect 321908 136368 324379 136370
rect 321908 136312 324318 136368
rect 324374 136312 324379 136368
rect 321908 136310 324379 136312
rect 324313 136307 324379 136310
rect 252461 136234 252527 136237
rect 248952 136232 252527 136234
rect 248952 136176 252466 136232
rect 252522 136176 252527 136232
rect 248952 136174 252527 136176
rect 252461 136171 252527 136174
rect 307569 136234 307635 136237
rect 307569 136232 310040 136234
rect 307569 136176 307574 136232
rect 307630 136176 310040 136232
rect 307569 136174 310040 136176
rect 307569 136171 307635 136174
rect 214741 136096 217242 136098
rect 214741 136040 214746 136096
rect 214802 136040 217242 136096
rect 214741 136038 217242 136040
rect 214741 136035 214807 136038
rect 213913 135690 213979 135693
rect 217182 135690 217242 135932
rect 252369 135690 252435 135693
rect 213913 135688 217242 135690
rect 213913 135632 213918 135688
rect 213974 135632 217242 135688
rect 213913 135630 217242 135632
rect 248952 135688 252435 135690
rect 248952 135632 252374 135688
rect 252430 135632 252435 135688
rect 248952 135630 252435 135632
rect 213913 135627 213979 135630
rect 252369 135627 252435 135630
rect 306741 135690 306807 135693
rect 306741 135688 310040 135690
rect 306741 135632 306746 135688
rect 306802 135632 310040 135688
rect 306741 135630 310040 135632
rect 306741 135627 306807 135630
rect 324497 135554 324563 135557
rect 321908 135552 324563 135554
rect 321908 135496 324502 135552
rect 324558 135496 324563 135552
rect 321908 135494 324563 135496
rect 324497 135491 324563 135494
rect 200070 135358 217242 135418
rect 169150 135220 169156 135284
rect 169220 135282 169226 135284
rect 200070 135282 200130 135358
rect 169220 135222 200130 135282
rect 217182 135252 217242 135358
rect 252277 135282 252343 135285
rect 248952 135280 252343 135282
rect 248952 135224 252282 135280
rect 252338 135224 252343 135280
rect 248952 135222 252343 135224
rect 169220 135220 169226 135222
rect 252277 135219 252343 135222
rect 307661 135282 307727 135285
rect 307661 135280 310040 135282
rect 307661 135224 307666 135280
rect 307722 135224 310040 135280
rect 307661 135222 310040 135224
rect 307661 135219 307727 135222
rect 308581 134874 308647 134877
rect 308581 134872 310040 134874
rect 308581 134816 308586 134872
rect 308642 134816 310040 134872
rect 308581 134814 310040 134816
rect 308581 134811 308647 134814
rect 252461 134738 252527 134741
rect 324313 134738 324379 134741
rect 248952 134736 252527 134738
rect 248952 134680 252466 134736
rect 252522 134680 252527 134736
rect 248952 134678 252527 134680
rect 321908 134736 324379 134738
rect 321908 134680 324318 134736
rect 324374 134680 324379 134736
rect 321908 134678 324379 134680
rect 252461 134675 252527 134678
rect 324313 134675 324379 134678
rect 166390 134132 166396 134196
rect 166460 134194 166466 134196
rect 217182 134194 217242 134572
rect 307661 134466 307727 134469
rect 307661 134464 310040 134466
rect 307661 134408 307666 134464
rect 307722 134408 310040 134464
rect 307661 134406 310040 134408
rect 307661 134403 307727 134406
rect 321502 134404 321508 134468
rect 321572 134404 321578 134468
rect 252369 134330 252435 134333
rect 248952 134328 252435 134330
rect 248952 134272 252374 134328
rect 252430 134272 252435 134328
rect 248952 134270 252435 134272
rect 252369 134267 252435 134270
rect 166460 134134 217242 134194
rect 166460 134132 166466 134134
rect 253054 134132 253060 134196
rect 253124 134194 253130 134196
rect 253124 134134 296730 134194
rect 253124 134132 253130 134134
rect 213913 134058 213979 134061
rect 296670 134058 296730 134134
rect 213913 134056 217242 134058
rect 213913 134000 213918 134056
rect 213974 134000 217242 134056
rect 213913 133998 217242 134000
rect 296670 133998 310040 134058
rect 321510 134028 321570 134404
rect 213913 133995 213979 133998
rect 217182 133892 217242 133998
rect 252461 133786 252527 133789
rect 248952 133784 252527 133786
rect 248952 133728 252466 133784
rect 252522 133728 252527 133784
rect 248952 133726 252527 133728
rect 252461 133723 252527 133726
rect 306557 133650 306623 133653
rect 306557 133648 310040 133650
rect 306557 133592 306562 133648
rect 306618 133592 310040 133648
rect 306557 133590 310040 133592
rect 306557 133587 306623 133590
rect 252369 133378 252435 133381
rect 248952 133376 252435 133378
rect 214005 132834 214071 132837
rect 217182 132834 217242 133348
rect 248952 133320 252374 133376
rect 252430 133320 252435 133376
rect 248952 133318 252435 133320
rect 252369 133315 252435 133318
rect 307109 133242 307175 133245
rect 324313 133242 324379 133245
rect 307109 133240 310040 133242
rect 307109 133184 307114 133240
rect 307170 133184 310040 133240
rect 307109 133182 310040 133184
rect 321908 133240 324379 133242
rect 321908 133184 324318 133240
rect 324374 133184 324379 133240
rect 321908 133182 324379 133184
rect 307109 133179 307175 133182
rect 324313 133179 324379 133182
rect 252277 132834 252343 132837
rect 214005 132832 217242 132834
rect 214005 132776 214010 132832
rect 214066 132776 217242 132832
rect 214005 132774 217242 132776
rect 248952 132832 252343 132834
rect 248952 132776 252282 132832
rect 252338 132776 252343 132832
rect 248952 132774 252343 132776
rect 214005 132771 214071 132774
rect 252277 132771 252343 132774
rect 307661 132698 307727 132701
rect 307661 132696 310040 132698
rect 213913 132562 213979 132565
rect 213913 132560 216874 132562
rect 213913 132504 213918 132560
rect 213974 132510 216874 132560
rect 217366 132510 217426 132668
rect 307661 132640 307666 132696
rect 307722 132640 310040 132696
rect 307661 132638 310040 132640
rect 307661 132635 307727 132638
rect 213974 132504 217426 132510
rect 213913 132502 217426 132504
rect 213913 132499 213979 132502
rect 216814 132450 217426 132502
rect 252461 132426 252527 132429
rect 324957 132426 325023 132429
rect 248952 132424 252527 132426
rect 248952 132368 252466 132424
rect 252522 132368 252527 132424
rect 248952 132366 252527 132368
rect 321908 132424 325023 132426
rect 321908 132368 324962 132424
rect 325018 132368 325023 132424
rect 321908 132366 325023 132368
rect 252461 132363 252527 132366
rect 324957 132363 325023 132366
rect 306557 132290 306623 132293
rect 306557 132288 310040 132290
rect 306557 132232 306562 132288
rect 306618 132232 310040 132288
rect 306557 132230 310040 132232
rect 306557 132227 306623 132230
rect 214005 131474 214071 131477
rect 217182 131474 217242 131988
rect 252369 131882 252435 131885
rect 248952 131880 252435 131882
rect 248952 131824 252374 131880
rect 252430 131824 252435 131880
rect 248952 131822 252435 131824
rect 252369 131819 252435 131822
rect 306925 131882 306991 131885
rect 306925 131880 310040 131882
rect 306925 131824 306930 131880
rect 306986 131824 310040 131880
rect 306925 131822 310040 131824
rect 306925 131819 306991 131822
rect 264513 131746 264579 131749
rect 307518 131746 307524 131748
rect 264513 131744 307524 131746
rect 264513 131688 264518 131744
rect 264574 131688 307524 131744
rect 264513 131686 307524 131688
rect 264513 131683 264579 131686
rect 307518 131684 307524 131686
rect 307588 131684 307594 131748
rect 327022 131746 327028 131748
rect 321908 131686 327028 131746
rect 327022 131684 327028 131686
rect 327092 131684 327098 131748
rect 252277 131474 252343 131477
rect 214005 131472 217242 131474
rect 214005 131416 214010 131472
rect 214066 131416 217242 131472
rect 214005 131414 217242 131416
rect 248952 131472 252343 131474
rect 248952 131416 252282 131472
rect 252338 131416 252343 131472
rect 248952 131414 252343 131416
rect 214005 131411 214071 131414
rect 252277 131411 252343 131414
rect 304206 131412 304212 131476
rect 304276 131474 304282 131476
rect 304276 131414 310040 131474
rect 304276 131412 304282 131414
rect 213913 131202 213979 131205
rect 213913 131200 216874 131202
rect 213913 131144 213918 131200
rect 213974 131144 216874 131200
rect 213913 131142 216874 131144
rect 213913 131139 213979 131142
rect 216814 131066 216874 131142
rect 217366 131066 217426 131308
rect 216814 131006 217426 131066
rect 307477 131066 307543 131069
rect 307477 131064 310040 131066
rect 307477 131008 307482 131064
rect 307538 131008 310040 131064
rect 307477 131006 310040 131008
rect 307477 131003 307543 131006
rect 252461 130930 252527 130933
rect 324313 130930 324379 130933
rect 248952 130928 252527 130930
rect 248952 130872 252466 130928
rect 252522 130872 252527 130928
rect 248952 130870 252527 130872
rect 321908 130928 324379 130930
rect 321908 130872 324318 130928
rect 324374 130872 324379 130928
rect 321908 130870 324379 130872
rect 252461 130867 252527 130870
rect 324313 130867 324379 130870
rect 166206 130052 166212 130116
rect 166276 130114 166282 130116
rect 217182 130114 217242 130628
rect 309550 130554 310132 130614
rect 252369 130522 252435 130525
rect 248952 130520 252435 130522
rect 248952 130464 252374 130520
rect 252430 130464 252435 130520
rect 248952 130462 252435 130464
rect 252369 130459 252435 130462
rect 252277 130114 252343 130117
rect 166276 130054 217242 130114
rect 248952 130112 252343 130114
rect 248952 130056 252282 130112
rect 252338 130056 252343 130112
rect 248952 130054 252343 130056
rect 166276 130052 166282 130054
rect 252277 130051 252343 130054
rect 305494 130052 305500 130116
rect 305564 130114 305570 130116
rect 309550 130114 309610 130554
rect 305564 130054 309610 130114
rect 309734 130146 310132 130206
rect 305564 130052 305570 130054
rect 307661 129978 307727 129981
rect 309734 129978 309794 130146
rect 324405 130114 324471 130117
rect 321908 130112 324471 130114
rect 321908 130056 324410 130112
rect 324466 130056 324471 130112
rect 321908 130054 324471 130056
rect 324405 130051 324471 130054
rect 307661 129976 309794 129978
rect 213913 129842 213979 129845
rect 213913 129840 216874 129842
rect 213913 129784 213918 129840
rect 213974 129784 216874 129840
rect 213913 129782 216874 129784
rect 213913 129779 213979 129782
rect 216814 129706 216874 129782
rect 217366 129706 217426 129948
rect 307661 129920 307666 129976
rect 307722 129920 309794 129976
rect 307661 129918 309794 129920
rect 307661 129915 307727 129918
rect 307293 129842 307359 129845
rect 307293 129840 310040 129842
rect 307293 129784 307298 129840
rect 307354 129784 310040 129840
rect 307293 129782 310040 129784
rect 307293 129779 307359 129782
rect 216814 129646 217426 129706
rect 252461 129570 252527 129573
rect 248952 129568 252527 129570
rect 248952 129512 252466 129568
rect 252522 129512 252527 129568
rect 248952 129510 252527 129512
rect 252461 129507 252527 129510
rect 324313 129434 324379 129437
rect 321908 129432 324379 129434
rect 321908 129376 324318 129432
rect 324374 129376 324379 129432
rect 321908 129374 324379 129376
rect 324313 129371 324379 129374
rect 66161 129298 66227 129301
rect 68142 129298 68816 129304
rect 66161 129296 68816 129298
rect 66161 129240 66166 129296
rect 66222 129244 68816 129296
rect 307569 129298 307635 129301
rect 307569 129296 310040 129298
rect 66222 129240 68202 129244
rect 66161 129238 68202 129240
rect 66161 129235 66227 129238
rect 213913 128890 213979 128893
rect 217182 128890 217242 129268
rect 307569 129240 307574 129296
rect 307630 129240 310040 129296
rect 307569 129238 310040 129240
rect 307569 129235 307635 129238
rect 252093 129162 252159 129165
rect 248952 129160 252159 129162
rect 248952 129104 252098 129160
rect 252154 129104 252159 129160
rect 248952 129102 252159 129104
rect 252093 129099 252159 129102
rect 213913 128888 217242 128890
rect 213913 128832 213918 128888
rect 213974 128832 217242 128888
rect 213913 128830 217242 128832
rect 307661 128890 307727 128893
rect 307661 128888 310040 128890
rect 307661 128832 307666 128888
rect 307722 128832 310040 128888
rect 307661 128830 310040 128832
rect 213913 128827 213979 128830
rect 307661 128827 307727 128830
rect 168966 128556 168972 128620
rect 169036 128618 169042 128620
rect 169036 128558 200130 128618
rect 169036 128556 169042 128558
rect 200070 128482 200130 128558
rect 217366 128482 217426 128724
rect 252369 128618 252435 128621
rect 324405 128618 324471 128621
rect 248952 128616 252435 128618
rect 248952 128560 252374 128616
rect 252430 128560 252435 128616
rect 248952 128558 252435 128560
rect 321908 128616 324471 128618
rect 321908 128560 324410 128616
rect 324466 128560 324471 128616
rect 321908 128558 324471 128560
rect 252369 128555 252435 128558
rect 324405 128555 324471 128558
rect 200070 128422 217426 128482
rect 307477 128482 307543 128485
rect 307477 128480 310040 128482
rect 307477 128424 307482 128480
rect 307538 128424 310040 128480
rect 307477 128422 310040 128424
rect 307477 128419 307543 128422
rect 252461 128210 252527 128213
rect 248952 128208 252527 128210
rect 248952 128152 252466 128208
rect 252522 128152 252527 128208
rect 248952 128150 252527 128152
rect 252461 128147 252527 128150
rect 67449 128074 67515 128077
rect 68142 128074 68816 128080
rect 67449 128072 68816 128074
rect 67449 128016 67454 128072
rect 67510 128020 68816 128072
rect 307477 128074 307543 128077
rect 307477 128072 310040 128074
rect 67510 128016 68202 128020
rect 67449 128014 68202 128016
rect 67449 128011 67515 128014
rect 217182 127530 217242 128044
rect 307477 128016 307482 128072
rect 307538 128016 310040 128072
rect 307477 128014 310040 128016
rect 307477 128011 307543 128014
rect 324313 127802 324379 127805
rect 321908 127800 324379 127802
rect 321908 127744 324318 127800
rect 324374 127744 324379 127800
rect 321908 127742 324379 127744
rect 324313 127739 324379 127742
rect 252277 127666 252343 127669
rect 248952 127664 252343 127666
rect 248952 127608 252282 127664
rect 252338 127608 252343 127664
rect 248952 127606 252343 127608
rect 252277 127603 252343 127606
rect 307569 127666 307635 127669
rect 307569 127664 310040 127666
rect 307569 127608 307574 127664
rect 307630 127608 310040 127664
rect 307569 127606 310040 127608
rect 307569 127603 307635 127606
rect 200070 127470 217242 127530
rect 321645 127530 321711 127533
rect 321645 127528 321754 127530
rect 321645 127472 321650 127528
rect 321706 127472 321754 127528
rect 168230 127060 168236 127124
rect 168300 127122 168306 127124
rect 200070 127122 200130 127470
rect 321645 127467 321754 127472
rect 168300 127062 200130 127122
rect 213913 127122 213979 127125
rect 217182 127122 217242 127364
rect 252369 127258 252435 127261
rect 248952 127256 252435 127258
rect 248952 127200 252374 127256
rect 252430 127200 252435 127256
rect 248952 127198 252435 127200
rect 252369 127195 252435 127198
rect 307661 127258 307727 127261
rect 307661 127256 310040 127258
rect 307661 127200 307666 127256
rect 307722 127200 310040 127256
rect 307661 127198 310040 127200
rect 307661 127195 307727 127198
rect 213913 127120 217242 127122
rect 213913 127064 213918 127120
rect 213974 127064 217242 127120
rect 321694 127092 321754 127467
rect 213913 127062 217242 127064
rect 168300 127060 168306 127062
rect 213913 127059 213979 127062
rect 306557 126850 306623 126853
rect 306557 126848 310040 126850
rect 306557 126792 306562 126848
rect 306618 126792 310040 126848
rect 306557 126790 310040 126792
rect 306557 126787 306623 126790
rect 252461 126714 252527 126717
rect 248952 126712 252527 126714
rect 65149 126306 65215 126309
rect 68142 126306 68816 126312
rect 65149 126304 68816 126306
rect 65149 126248 65154 126304
rect 65210 126252 68816 126304
rect 65210 126248 68202 126252
rect 65149 126246 68202 126248
rect 65149 126243 65215 126246
rect 214005 126170 214071 126173
rect 217182 126170 217242 126684
rect 248952 126656 252466 126712
rect 252522 126656 252527 126712
rect 248952 126654 252527 126656
rect 252461 126651 252527 126654
rect 306966 126380 306972 126444
rect 307036 126442 307042 126444
rect 307036 126382 310040 126442
rect 307036 126380 307042 126382
rect 252185 126306 252251 126309
rect 324497 126306 324563 126309
rect 248952 126304 252251 126306
rect 248952 126248 252190 126304
rect 252246 126248 252251 126304
rect 248952 126246 252251 126248
rect 321908 126304 324563 126306
rect 321908 126248 324502 126304
rect 324558 126248 324563 126304
rect 321908 126246 324563 126248
rect 252185 126243 252251 126246
rect 324497 126243 324563 126246
rect 214005 126168 217242 126170
rect 214005 126112 214010 126168
rect 214066 126112 217242 126168
rect 214005 126110 217242 126112
rect 214005 126107 214071 126110
rect 582925 126034 582991 126037
rect 583520 126034 584960 126124
rect 582925 126032 584960 126034
rect 213913 125762 213979 125765
rect 217182 125762 217242 126004
rect 582925 125976 582930 126032
rect 582986 125976 584960 126032
rect 582925 125974 584960 125976
rect 582925 125971 582991 125974
rect 307661 125898 307727 125901
rect 307661 125896 310040 125898
rect 307661 125840 307666 125896
rect 307722 125840 310040 125896
rect 583520 125884 584960 125974
rect 307661 125838 310040 125840
rect 307661 125835 307727 125838
rect 251725 125762 251791 125765
rect 213913 125760 217242 125762
rect 213913 125704 213918 125760
rect 213974 125704 217242 125760
rect 213913 125702 217242 125704
rect 248952 125760 251791 125762
rect 248952 125704 251730 125760
rect 251786 125704 251791 125760
rect 248952 125702 251791 125704
rect 213913 125699 213979 125702
rect 251725 125699 251791 125702
rect 306557 125490 306623 125493
rect 324313 125490 324379 125493
rect 306557 125488 310040 125490
rect 306557 125432 306562 125488
rect 306618 125432 310040 125488
rect 306557 125430 310040 125432
rect 321908 125488 324379 125490
rect 321908 125432 324318 125488
rect 324374 125432 324379 125488
rect 321908 125430 324379 125432
rect 306557 125427 306623 125430
rect 324313 125427 324379 125430
rect 252277 125354 252343 125357
rect 248952 125352 252343 125354
rect 65517 125218 65583 125221
rect 68142 125218 68816 125224
rect 65517 125216 68816 125218
rect 65517 125160 65522 125216
rect 65578 125164 68816 125216
rect 65578 125160 68202 125164
rect 65517 125158 68202 125160
rect 65517 125155 65583 125158
rect 214005 124810 214071 124813
rect 217182 124810 217242 125324
rect 248952 125296 252282 125352
rect 252338 125296 252343 125352
rect 248952 125294 252343 125296
rect 252277 125291 252343 125294
rect 307569 125082 307635 125085
rect 307569 125080 310040 125082
rect 307569 125024 307574 125080
rect 307630 125024 310040 125080
rect 307569 125022 310040 125024
rect 307569 125019 307635 125022
rect 252461 124810 252527 124813
rect 214005 124808 217242 124810
rect 214005 124752 214010 124808
rect 214066 124752 217242 124808
rect 214005 124750 217242 124752
rect 248952 124808 252527 124810
rect 248952 124752 252466 124808
rect 252522 124752 252527 124808
rect 248952 124750 252527 124752
rect 214005 124747 214071 124750
rect 252461 124747 252527 124750
rect 307661 124674 307727 124677
rect 307661 124672 310040 124674
rect 213913 124402 213979 124405
rect 217182 124402 217242 124644
rect 307661 124616 307666 124672
rect 307722 124616 310040 124672
rect 307661 124614 310040 124616
rect 307661 124611 307727 124614
rect 252369 124402 252435 124405
rect 213913 124400 217242 124402
rect 213913 124344 213918 124400
rect 213974 124344 217242 124400
rect 213913 124342 217242 124344
rect 248952 124400 252435 124402
rect 248952 124344 252374 124400
rect 252430 124344 252435 124400
rect 248952 124342 252435 124344
rect 213913 124339 213979 124342
rect 252369 124339 252435 124342
rect 307477 124266 307543 124269
rect 321878 124266 321938 124780
rect 339718 124266 339724 124268
rect 307477 124264 310040 124266
rect 307477 124208 307482 124264
rect 307538 124208 310040 124264
rect 307477 124206 310040 124208
rect 321878 124206 339724 124266
rect 307477 124203 307543 124206
rect 339718 124204 339724 124206
rect 339788 124204 339794 124268
rect -960 123572 480 123812
rect 66069 123586 66135 123589
rect 68142 123586 68816 123592
rect 66069 123584 68816 123586
rect 66069 123528 66074 123584
rect 66130 123532 68816 123584
rect 214005 123586 214071 123589
rect 217182 123586 217242 124100
rect 252461 123994 252527 123997
rect 324313 123994 324379 123997
rect 248952 123992 252527 123994
rect 248952 123936 252466 123992
rect 252522 123936 252527 123992
rect 248952 123934 252527 123936
rect 321908 123992 324379 123994
rect 321908 123936 324318 123992
rect 324374 123936 324379 123992
rect 321908 123934 324379 123936
rect 252461 123931 252527 123934
rect 324313 123931 324379 123934
rect 307477 123858 307543 123861
rect 307477 123856 310040 123858
rect 307477 123800 307482 123856
rect 307538 123800 310040 123856
rect 307477 123798 310040 123800
rect 307477 123795 307543 123798
rect 214005 123584 217242 123586
rect 66130 123528 68202 123532
rect 66069 123526 68202 123528
rect 214005 123528 214010 123584
rect 214066 123528 217242 123584
rect 214005 123526 217242 123528
rect 66069 123523 66135 123526
rect 214005 123523 214071 123526
rect 252369 123450 252435 123453
rect 248952 123448 252435 123450
rect 213913 123178 213979 123181
rect 217182 123178 217242 123420
rect 248952 123392 252374 123448
rect 252430 123392 252435 123448
rect 248952 123390 252435 123392
rect 252369 123387 252435 123390
rect 307569 123450 307635 123453
rect 307569 123448 310040 123450
rect 307569 123392 307574 123448
rect 307630 123392 310040 123448
rect 307569 123390 310040 123392
rect 307569 123387 307635 123390
rect 324405 123178 324471 123181
rect 213913 123176 217242 123178
rect 213913 123120 213918 123176
rect 213974 123120 217242 123176
rect 213913 123118 217242 123120
rect 321908 123176 324471 123178
rect 321908 123120 324410 123176
rect 324466 123120 324471 123176
rect 321908 123118 324471 123120
rect 213913 123115 213979 123118
rect 324405 123115 324471 123118
rect 252277 123042 252343 123045
rect 248952 123040 252343 123042
rect 248952 122984 252282 123040
rect 252338 122984 252343 123040
rect 248952 122982 252343 122984
rect 252277 122979 252343 122982
rect 307661 123042 307727 123045
rect 307661 123040 310040 123042
rect 307661 122984 307666 123040
rect 307722 122984 310040 123040
rect 307661 122982 310040 122984
rect 307661 122979 307727 122982
rect 67357 122634 67423 122637
rect 68142 122634 68816 122640
rect 67357 122632 68816 122634
rect 67357 122576 67362 122632
rect 67418 122580 68816 122632
rect 67418 122576 68202 122580
rect 67357 122574 68202 122576
rect 67357 122571 67423 122574
rect 214005 122226 214071 122229
rect 217182 122226 217242 122740
rect 252461 122498 252527 122501
rect 248952 122496 252527 122498
rect 248952 122440 252466 122496
rect 252522 122440 252527 122496
rect 248952 122438 252527 122440
rect 252461 122435 252527 122438
rect 307569 122498 307635 122501
rect 324313 122498 324379 122501
rect 307569 122496 310040 122498
rect 307569 122440 307574 122496
rect 307630 122440 310040 122496
rect 307569 122438 310040 122440
rect 321908 122496 324379 122498
rect 321908 122440 324318 122496
rect 324374 122440 324379 122496
rect 321908 122438 324379 122440
rect 307569 122435 307635 122438
rect 324313 122435 324379 122438
rect 214005 122224 217242 122226
rect 214005 122168 214010 122224
rect 214066 122168 217242 122224
rect 214005 122166 217242 122168
rect 214005 122163 214071 122166
rect 252277 122090 252343 122093
rect 248952 122088 252343 122090
rect 213913 121546 213979 121549
rect 217182 121546 217242 122060
rect 248952 122032 252282 122088
rect 252338 122032 252343 122088
rect 248952 122030 252343 122032
rect 252277 122027 252343 122030
rect 307661 122090 307727 122093
rect 307661 122088 310040 122090
rect 307661 122032 307666 122088
rect 307722 122032 310040 122088
rect 307661 122030 310040 122032
rect 307661 122027 307727 122030
rect 307477 121682 307543 121685
rect 323025 121682 323091 121685
rect 307477 121680 310040 121682
rect 307477 121624 307482 121680
rect 307538 121624 310040 121680
rect 307477 121622 310040 121624
rect 321908 121680 323091 121682
rect 321908 121624 323030 121680
rect 323086 121624 323091 121680
rect 321908 121622 323091 121624
rect 307477 121619 307543 121622
rect 323025 121619 323091 121622
rect 252369 121546 252435 121549
rect 213913 121544 217242 121546
rect 213913 121488 213918 121544
rect 213974 121488 217242 121544
rect 213913 121486 217242 121488
rect 248952 121544 252435 121546
rect 248952 121488 252374 121544
rect 252430 121488 252435 121544
rect 248952 121486 252435 121488
rect 213913 121483 213979 121486
rect 252369 121483 252435 121486
rect 67541 120866 67607 120869
rect 68142 120866 68816 120872
rect 67541 120864 68816 120866
rect 67541 120808 67546 120864
rect 67602 120812 68816 120864
rect 214005 120866 214071 120869
rect 217182 120866 217242 121380
rect 307109 121274 307175 121277
rect 307109 121272 310040 121274
rect 307109 121216 307114 121272
rect 307170 121216 310040 121272
rect 307109 121214 310040 121216
rect 307109 121211 307175 121214
rect 252461 121138 252527 121141
rect 248952 121136 252527 121138
rect 248952 121080 252466 121136
rect 252522 121080 252527 121136
rect 248952 121078 252527 121080
rect 252461 121075 252527 121078
rect 214005 120864 217242 120866
rect 67602 120808 68202 120812
rect 67541 120806 68202 120808
rect 214005 120808 214010 120864
rect 214066 120808 217242 120864
rect 214005 120806 217242 120808
rect 307569 120866 307635 120869
rect 322933 120866 322999 120869
rect 307569 120864 310040 120866
rect 307569 120808 307574 120864
rect 307630 120808 310040 120864
rect 307569 120806 310040 120808
rect 321908 120864 322999 120866
rect 321908 120808 322938 120864
rect 322994 120808 322999 120864
rect 321908 120806 322999 120808
rect 67541 120803 67607 120806
rect 214005 120803 214071 120806
rect 307569 120803 307635 120806
rect 322933 120803 322999 120806
rect 213913 120458 213979 120461
rect 217182 120458 217242 120700
rect 252369 120594 252435 120597
rect 248952 120592 252435 120594
rect 248952 120536 252374 120592
rect 252430 120536 252435 120592
rect 248952 120534 252435 120536
rect 252369 120531 252435 120534
rect 213913 120456 217242 120458
rect 213913 120400 213918 120456
rect 213974 120400 217242 120456
rect 213913 120398 217242 120400
rect 307661 120458 307727 120461
rect 307661 120456 310040 120458
rect 307661 120400 307666 120456
rect 307722 120400 310040 120456
rect 307661 120398 310040 120400
rect 213913 120395 213979 120398
rect 307661 120395 307727 120398
rect 252461 120186 252527 120189
rect 324313 120186 324379 120189
rect 248952 120184 252527 120186
rect 248952 120128 252466 120184
rect 252522 120128 252527 120184
rect 248952 120126 252527 120128
rect 321908 120184 324379 120186
rect 321908 120128 324318 120184
rect 324374 120128 324379 120184
rect 321908 120126 324379 120128
rect 252461 120123 252527 120126
rect 324313 120123 324379 120126
rect 307109 120050 307175 120053
rect 307109 120048 310040 120050
rect 213361 119642 213427 119645
rect 217182 119642 217242 120020
rect 307109 119992 307114 120048
rect 307170 119992 310040 120048
rect 307109 119990 310040 119992
rect 307109 119987 307175 119990
rect 321553 119914 321619 119917
rect 321510 119912 321619 119914
rect 321510 119856 321558 119912
rect 321614 119856 321619 119912
rect 321510 119851 321619 119856
rect 252461 119642 252527 119645
rect 213361 119640 217242 119642
rect 213361 119584 213366 119640
rect 213422 119584 217242 119640
rect 213361 119582 217242 119584
rect 248952 119640 252527 119642
rect 248952 119584 252466 119640
rect 252522 119584 252527 119640
rect 248952 119582 252527 119584
rect 213361 119579 213427 119582
rect 252461 119579 252527 119582
rect 307569 119642 307635 119645
rect 307569 119640 310040 119642
rect 307569 119584 307574 119640
rect 307630 119584 310040 119640
rect 307569 119582 310040 119584
rect 307569 119579 307635 119582
rect 214005 119098 214071 119101
rect 217182 119098 217242 119476
rect 321510 119340 321570 119851
rect 252277 119234 252343 119237
rect 248952 119232 252343 119234
rect 248952 119176 252282 119232
rect 252338 119176 252343 119232
rect 248952 119174 252343 119176
rect 252277 119171 252343 119174
rect 214005 119096 217242 119098
rect 214005 119040 214010 119096
rect 214066 119040 217242 119096
rect 214005 119038 217242 119040
rect 307661 119098 307727 119101
rect 307661 119096 310040 119098
rect 307661 119040 307666 119096
rect 307722 119040 310040 119096
rect 307661 119038 310040 119040
rect 214005 119035 214071 119038
rect 307661 119035 307727 119038
rect 213913 118962 213979 118965
rect 213913 118960 217242 118962
rect 213913 118904 213918 118960
rect 213974 118904 217242 118960
rect 213913 118902 217242 118904
rect 213913 118899 213979 118902
rect 217182 118796 217242 118902
rect 252001 118826 252067 118829
rect 248952 118824 252067 118826
rect 248952 118768 252006 118824
rect 252062 118768 252067 118824
rect 248952 118766 252067 118768
rect 252001 118763 252067 118766
rect 306557 118690 306623 118693
rect 306557 118688 310040 118690
rect 306557 118632 306562 118688
rect 306618 118632 310040 118688
rect 306557 118630 310040 118632
rect 306557 118627 306623 118630
rect 324313 118554 324379 118557
rect 321908 118552 324379 118554
rect 321908 118496 324318 118552
rect 324374 118496 324379 118552
rect 321908 118494 324379 118496
rect 324313 118491 324379 118494
rect 252461 118282 252527 118285
rect 248952 118280 252527 118282
rect 248952 118224 252466 118280
rect 252522 118224 252527 118280
rect 248952 118222 252527 118224
rect 252461 118219 252527 118222
rect 307569 118282 307635 118285
rect 307569 118280 310040 118282
rect 307569 118224 307574 118280
rect 307630 118224 310040 118280
rect 307569 118222 310040 118224
rect 307569 118219 307635 118222
rect 214005 117602 214071 117605
rect 217182 117602 217242 118116
rect 252461 117874 252527 117877
rect 248952 117872 252527 117874
rect 248952 117816 252466 117872
rect 252522 117816 252527 117872
rect 248952 117814 252527 117816
rect 252461 117811 252527 117814
rect 307661 117874 307727 117877
rect 324405 117874 324471 117877
rect 307661 117872 310040 117874
rect 307661 117816 307666 117872
rect 307722 117816 310040 117872
rect 307661 117814 310040 117816
rect 321908 117872 324471 117874
rect 321908 117816 324410 117872
rect 324466 117816 324471 117872
rect 321908 117814 324471 117816
rect 307661 117811 307727 117814
rect 324405 117811 324471 117814
rect 214005 117600 217242 117602
rect 214005 117544 214010 117600
rect 214066 117544 217242 117600
rect 214005 117542 217242 117544
rect 214005 117539 214071 117542
rect 307109 117466 307175 117469
rect 307109 117464 310040 117466
rect 213913 117330 213979 117333
rect 213913 117328 216874 117330
rect 213913 117272 213918 117328
rect 213974 117272 216874 117328
rect 213913 117270 216874 117272
rect 213913 117267 213979 117270
rect 216814 117194 216874 117270
rect 217366 117194 217426 117436
rect 307109 117408 307114 117464
rect 307170 117408 310040 117464
rect 307109 117406 310040 117408
rect 307109 117403 307175 117406
rect 252369 117330 252435 117333
rect 248952 117328 252435 117330
rect 248952 117272 252374 117328
rect 252430 117272 252435 117328
rect 248952 117270 252435 117272
rect 252369 117267 252435 117270
rect 216814 117134 217426 117194
rect 307661 117058 307727 117061
rect 307661 117056 310040 117058
rect 307661 117000 307666 117056
rect 307722 117000 310040 117056
rect 307661 116998 310040 117000
rect 307661 116995 307727 116998
rect 252461 116922 252527 116925
rect 248952 116920 252527 116922
rect 248952 116864 252466 116920
rect 252522 116864 252527 116920
rect 248952 116862 252527 116864
rect 252461 116859 252527 116862
rect 214005 116242 214071 116245
rect 217182 116242 217242 116756
rect 306925 116650 306991 116653
rect 306925 116648 310040 116650
rect 306925 116592 306930 116648
rect 306986 116592 310040 116648
rect 306925 116590 310040 116592
rect 306925 116587 306991 116590
rect 321878 116514 321938 117028
rect 321878 116454 325710 116514
rect 252369 116378 252435 116381
rect 324313 116378 324379 116381
rect 248952 116376 252435 116378
rect 248952 116320 252374 116376
rect 252430 116320 252435 116376
rect 248952 116318 252435 116320
rect 321908 116376 324379 116378
rect 321908 116320 324318 116376
rect 324374 116320 324379 116376
rect 321908 116318 324379 116320
rect 252369 116315 252435 116318
rect 324313 116315 324379 116318
rect 214005 116240 217242 116242
rect 214005 116184 214010 116240
rect 214066 116184 217242 116240
rect 214005 116182 217242 116184
rect 307017 116242 307083 116245
rect 307017 116240 310040 116242
rect 307017 116184 307022 116240
rect 307078 116184 310040 116240
rect 307017 116182 310040 116184
rect 214005 116179 214071 116182
rect 307017 116179 307083 116182
rect 213913 115970 213979 115973
rect 213913 115968 216874 115970
rect 213913 115912 213918 115968
rect 213974 115912 216874 115968
rect 213913 115910 216874 115912
rect 213913 115907 213979 115910
rect 216814 115834 216874 115910
rect 217366 115834 217426 116076
rect 252461 115970 252527 115973
rect 248952 115968 252527 115970
rect 248952 115912 252466 115968
rect 252522 115912 252527 115968
rect 248952 115910 252527 115912
rect 325650 115970 325710 116454
rect 336774 115970 336780 115972
rect 325650 115910 336780 115970
rect 252461 115907 252527 115910
rect 336774 115908 336780 115910
rect 336844 115908 336850 115972
rect 216814 115774 217426 115834
rect 307109 115698 307175 115701
rect 307109 115696 310040 115698
rect 307109 115640 307114 115696
rect 307170 115640 310040 115696
rect 307109 115638 310040 115640
rect 307109 115635 307175 115638
rect 324313 115562 324379 115565
rect 321908 115560 324379 115562
rect 321908 115504 324318 115560
rect 324374 115504 324379 115560
rect 321908 115502 324379 115504
rect 324313 115499 324379 115502
rect 251817 115426 251883 115429
rect 248952 115424 251883 115426
rect 170254 115092 170260 115156
rect 170324 115154 170330 115156
rect 199377 115154 199443 115157
rect 170324 115152 199443 115154
rect 170324 115096 199382 115152
rect 199438 115096 199443 115152
rect 170324 115094 199443 115096
rect 170324 115092 170330 115094
rect 199377 115091 199443 115094
rect 213913 115018 213979 115021
rect 217182 115018 217242 115396
rect 248952 115368 251822 115424
rect 251878 115368 251883 115424
rect 248952 115366 251883 115368
rect 251817 115363 251883 115366
rect 307569 115290 307635 115293
rect 307569 115288 310040 115290
rect 307569 115232 307574 115288
rect 307630 115232 310040 115288
rect 307569 115230 310040 115232
rect 307569 115227 307635 115230
rect 252369 115018 252435 115021
rect 213913 115016 217242 115018
rect 213913 114960 213918 115016
rect 213974 114960 217242 115016
rect 213913 114958 217242 114960
rect 248952 115016 252435 115018
rect 248952 114960 252374 115016
rect 252430 114960 252435 115016
rect 248952 114958 252435 114960
rect 213913 114955 213979 114958
rect 252369 114955 252435 114958
rect 307661 114882 307727 114885
rect 307661 114880 310040 114882
rect 215017 114610 215083 114613
rect 217182 114610 217242 114852
rect 307661 114824 307666 114880
rect 307722 114824 310040 114880
rect 307661 114822 310040 114824
rect 307661 114819 307727 114822
rect 324405 114746 324471 114749
rect 321908 114744 324471 114746
rect 321908 114688 324410 114744
rect 324466 114688 324471 114744
rect 321908 114686 324471 114688
rect 324405 114683 324471 114686
rect 215017 114608 217242 114610
rect 215017 114552 215022 114608
rect 215078 114552 217242 114608
rect 215017 114550 217242 114552
rect 215017 114547 215083 114550
rect 251909 114474 251975 114477
rect 248952 114472 251975 114474
rect 248952 114416 251914 114472
rect 251970 114416 251975 114472
rect 248952 114414 251975 114416
rect 251909 114411 251975 114414
rect 307477 114474 307543 114477
rect 307477 114472 310040 114474
rect 307477 114416 307482 114472
rect 307538 114416 310040 114472
rect 307477 114414 310040 114416
rect 307477 114411 307543 114414
rect 213913 113658 213979 113661
rect 217182 113658 217242 114172
rect 252461 114066 252527 114069
rect 324313 114066 324379 114069
rect 248952 114064 252527 114066
rect 248952 114008 252466 114064
rect 252522 114008 252527 114064
rect 321908 114064 324379 114066
rect 248952 114006 252527 114008
rect 252461 114003 252527 114006
rect 309550 113962 310132 114022
rect 321908 114008 324318 114064
rect 324374 114008 324379 114064
rect 321908 114006 324379 114008
rect 324313 114003 324379 114006
rect 299974 113868 299980 113932
rect 300044 113930 300050 113932
rect 309550 113930 309610 113962
rect 300044 113870 309610 113930
rect 300044 113868 300050 113870
rect 213913 113656 217242 113658
rect 213913 113600 213918 113656
rect 213974 113600 217242 113656
rect 213913 113598 217242 113600
rect 307569 113658 307635 113661
rect 307569 113656 310040 113658
rect 307569 113600 307574 113656
rect 307630 113600 310040 113656
rect 307569 113598 310040 113600
rect 213913 113595 213979 113598
rect 307569 113595 307635 113598
rect 251725 113522 251791 113525
rect 248952 113520 251791 113522
rect 213453 113250 213519 113253
rect 217366 113250 217426 113492
rect 248952 113464 251730 113520
rect 251786 113464 251791 113520
rect 248952 113462 251791 113464
rect 251725 113459 251791 113462
rect 213453 113248 217426 113250
rect 213453 113192 213458 113248
rect 213514 113192 217426 113248
rect 213453 113190 217426 113192
rect 307661 113250 307727 113253
rect 324405 113250 324471 113253
rect 307661 113248 310040 113250
rect 307661 113192 307666 113248
rect 307722 113192 310040 113248
rect 307661 113190 310040 113192
rect 321908 113248 324471 113250
rect 321908 113192 324410 113248
rect 324466 113192 324471 113248
rect 321908 113190 324471 113192
rect 213453 113187 213519 113190
rect 307661 113187 307727 113190
rect 324405 113187 324471 113190
rect 252461 113114 252527 113117
rect 248952 113112 252527 113114
rect 248952 113056 252466 113112
rect 252522 113056 252527 113112
rect 248952 113054 252527 113056
rect 252461 113051 252527 113054
rect 582557 112842 582623 112845
rect 583520 112842 584960 112932
rect 582557 112840 584960 112842
rect 214005 112298 214071 112301
rect 217182 112298 217242 112812
rect 582557 112784 582562 112840
rect 582618 112784 584960 112840
rect 582557 112782 584960 112784
rect 582557 112779 582623 112782
rect 252369 112706 252435 112709
rect 248952 112704 252435 112706
rect 248952 112648 252374 112704
rect 252430 112648 252435 112704
rect 248952 112646 252435 112648
rect 252369 112643 252435 112646
rect 307661 112706 307727 112709
rect 307661 112704 310040 112706
rect 307661 112648 307666 112704
rect 307722 112648 310040 112704
rect 583520 112692 584960 112782
rect 307661 112646 310040 112648
rect 307661 112643 307727 112646
rect 324313 112434 324379 112437
rect 321908 112432 324379 112434
rect 321908 112376 324318 112432
rect 324374 112376 324379 112432
rect 321908 112374 324379 112376
rect 324313 112371 324379 112374
rect 214005 112296 217242 112298
rect 214005 112240 214010 112296
rect 214066 112240 217242 112296
rect 214005 112238 217242 112240
rect 307569 112298 307635 112301
rect 307569 112296 310040 112298
rect 307569 112240 307574 112296
rect 307630 112240 310040 112296
rect 307569 112238 310040 112240
rect 214005 112235 214071 112238
rect 307569 112235 307635 112238
rect 252461 112162 252527 112165
rect 248952 112160 252527 112162
rect 213913 111890 213979 111893
rect 217182 111890 217242 112132
rect 248952 112104 252466 112160
rect 252522 112104 252527 112160
rect 248952 112102 252527 112104
rect 252461 112099 252527 112102
rect 213913 111888 217242 111890
rect 213913 111832 213918 111888
rect 213974 111832 217242 111888
rect 213913 111830 217242 111832
rect 307661 111890 307727 111893
rect 307661 111888 310040 111890
rect 307661 111832 307666 111888
rect 307722 111832 310040 111888
rect 307661 111830 310040 111832
rect 213913 111827 213979 111830
rect 307661 111827 307727 111830
rect 168281 111754 168347 111757
rect 252461 111754 252527 111757
rect 164694 111752 168347 111754
rect 164694 111696 168286 111752
rect 168342 111696 168347 111752
rect 164694 111694 168347 111696
rect 248952 111752 252527 111754
rect 248952 111696 252466 111752
rect 252522 111696 252527 111752
rect 248952 111694 252527 111696
rect 168281 111691 168347 111694
rect 252461 111691 252527 111694
rect 307569 111482 307635 111485
rect 307569 111480 310040 111482
rect 214005 110938 214071 110941
rect 217182 110938 217242 111452
rect 307569 111424 307574 111480
rect 307630 111424 310040 111480
rect 307569 111422 310040 111424
rect 307569 111419 307635 111422
rect 252277 111210 252343 111213
rect 248952 111208 252343 111210
rect 248952 111152 252282 111208
rect 252338 111152 252343 111208
rect 248952 111150 252343 111152
rect 252277 111147 252343 111150
rect 307477 111074 307543 111077
rect 321878 111074 321938 111724
rect 331438 111074 331444 111076
rect 307477 111072 310040 111074
rect 307477 111016 307482 111072
rect 307538 111016 310040 111072
rect 307477 111014 310040 111016
rect 321878 111014 331444 111074
rect 307477 111011 307543 111014
rect 331438 111012 331444 111014
rect 331508 111012 331514 111076
rect 324313 110938 324379 110941
rect 214005 110936 217242 110938
rect 214005 110880 214010 110936
rect 214066 110880 217242 110936
rect 214005 110878 217242 110880
rect 321908 110936 324379 110938
rect 321908 110880 324318 110936
rect 324374 110880 324379 110936
rect 321908 110878 324379 110880
rect 214005 110875 214071 110878
rect 324313 110875 324379 110878
rect 252369 110802 252435 110805
rect 248952 110800 252435 110802
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 213913 110530 213979 110533
rect 217366 110530 217426 110772
rect 248952 110744 252374 110800
rect 252430 110744 252435 110800
rect 248952 110742 252435 110744
rect 252369 110739 252435 110742
rect 307661 110666 307727 110669
rect 307661 110664 310040 110666
rect 307661 110608 307666 110664
rect 307722 110608 310040 110664
rect 307661 110606 310040 110608
rect 307661 110603 307727 110606
rect 213913 110528 217426 110530
rect 213913 110472 213918 110528
rect 213974 110472 217426 110528
rect 213913 110470 217426 110472
rect 213913 110467 213979 110470
rect 252461 110258 252527 110261
rect 248952 110256 252527 110258
rect 167821 110122 167887 110125
rect 164694 110120 167887 110122
rect 164694 110064 167826 110120
rect 167882 110064 167887 110120
rect 164694 110062 167887 110064
rect 167821 110059 167887 110062
rect 214005 109714 214071 109717
rect 217182 109714 217242 110228
rect 248952 110200 252466 110256
rect 252522 110200 252527 110256
rect 248952 110198 252527 110200
rect 252461 110195 252527 110198
rect 307477 110258 307543 110261
rect 307477 110256 310040 110258
rect 307477 110200 307482 110256
rect 307538 110200 310040 110256
rect 307477 110198 310040 110200
rect 307477 110195 307543 110198
rect 324313 110122 324379 110125
rect 321908 110120 324379 110122
rect 321908 110064 324318 110120
rect 324374 110064 324379 110120
rect 321908 110062 324379 110064
rect 324313 110059 324379 110062
rect 252369 109850 252435 109853
rect 248952 109848 252435 109850
rect 248952 109792 252374 109848
rect 252430 109792 252435 109848
rect 248952 109790 252435 109792
rect 252369 109787 252435 109790
rect 307569 109850 307635 109853
rect 307569 109848 310040 109850
rect 307569 109792 307574 109848
rect 307630 109792 310040 109848
rect 307569 109790 310040 109792
rect 307569 109787 307635 109790
rect 214005 109712 217242 109714
rect 214005 109656 214010 109712
rect 214066 109656 217242 109712
rect 214005 109654 217242 109656
rect 214005 109651 214071 109654
rect 213913 109306 213979 109309
rect 217182 109306 217242 109548
rect 324405 109442 324471 109445
rect 321908 109440 324471 109442
rect 321908 109384 324410 109440
rect 324466 109384 324471 109440
rect 321908 109382 324471 109384
rect 324405 109379 324471 109382
rect 252277 109306 252343 109309
rect 213913 109304 217242 109306
rect 213913 109248 213918 109304
rect 213974 109248 217242 109304
rect 213913 109246 217242 109248
rect 248952 109304 252343 109306
rect 248952 109248 252282 109304
rect 252338 109248 252343 109304
rect 248952 109246 252343 109248
rect 213913 109243 213979 109246
rect 252277 109243 252343 109246
rect 307661 109306 307727 109309
rect 307661 109304 310040 109306
rect 307661 109248 307666 109304
rect 307722 109248 310040 109304
rect 307661 109246 310040 109248
rect 307661 109243 307727 109246
rect 252461 108898 252527 108901
rect 248952 108896 252527 108898
rect 168097 108762 168163 108765
rect 164694 108760 168163 108762
rect 164694 108704 168102 108760
rect 168158 108704 168163 108760
rect 164694 108702 168163 108704
rect 168097 108699 168163 108702
rect 214649 108354 214715 108357
rect 217182 108354 217242 108868
rect 248952 108840 252466 108896
rect 252522 108840 252527 108896
rect 248952 108838 252527 108840
rect 252461 108835 252527 108838
rect 307661 108898 307727 108901
rect 307661 108896 310040 108898
rect 307661 108840 307666 108896
rect 307722 108840 310040 108896
rect 307661 108838 310040 108840
rect 307661 108835 307727 108838
rect 324405 108626 324471 108629
rect 321908 108624 324471 108626
rect 321908 108568 324410 108624
rect 324466 108568 324471 108624
rect 321908 108566 324471 108568
rect 324405 108563 324471 108566
rect 307569 108490 307635 108493
rect 307569 108488 310040 108490
rect 307569 108432 307574 108488
rect 307630 108432 310040 108488
rect 307569 108430 310040 108432
rect 307569 108427 307635 108430
rect 251725 108354 251791 108357
rect 214649 108352 217242 108354
rect 214649 108296 214654 108352
rect 214710 108296 217242 108352
rect 214649 108294 217242 108296
rect 248952 108352 251791 108354
rect 248952 108296 251730 108352
rect 251786 108296 251791 108352
rect 248952 108294 251791 108296
rect 214649 108291 214715 108294
rect 251725 108291 251791 108294
rect 213913 107946 213979 107949
rect 217182 107946 217242 108188
rect 305821 108082 305887 108085
rect 305821 108080 310040 108082
rect 305821 108024 305826 108080
rect 305882 108024 310040 108080
rect 305821 108022 310040 108024
rect 305821 108019 305887 108022
rect 252369 107946 252435 107949
rect 213913 107944 217242 107946
rect 213913 107888 213918 107944
rect 213974 107888 217242 107944
rect 213913 107886 217242 107888
rect 248952 107944 252435 107946
rect 248952 107888 252374 107944
rect 252430 107888 252435 107944
rect 248952 107886 252435 107888
rect 213913 107883 213979 107886
rect 252369 107883 252435 107886
rect 324313 107810 324379 107813
rect 321908 107808 324379 107810
rect 321908 107752 324318 107808
rect 324374 107752 324379 107808
rect 321908 107750 324379 107752
rect 324313 107747 324379 107750
rect 307477 107674 307543 107677
rect 307477 107672 310040 107674
rect 307477 107616 307482 107672
rect 307538 107616 310040 107672
rect 307477 107614 310040 107616
rect 307477 107611 307543 107614
rect 252461 107538 252527 107541
rect 248952 107536 252527 107538
rect 214005 106994 214071 106997
rect 217182 106994 217242 107508
rect 248952 107480 252466 107536
rect 252522 107480 252527 107536
rect 248952 107478 252527 107480
rect 252461 107475 252527 107478
rect 307661 107266 307727 107269
rect 307661 107264 310040 107266
rect 307661 107208 307666 107264
rect 307722 107208 310040 107264
rect 307661 107206 310040 107208
rect 307661 107203 307727 107206
rect 322974 107130 322980 107132
rect 321908 107070 322980 107130
rect 322974 107068 322980 107070
rect 323044 107068 323050 107132
rect 252277 106994 252343 106997
rect 214005 106992 217242 106994
rect 214005 106936 214010 106992
rect 214066 106936 217242 106992
rect 214005 106934 217242 106936
rect 248952 106992 252343 106994
rect 248952 106936 252282 106992
rect 252338 106936 252343 106992
rect 248952 106934 252343 106936
rect 214005 106931 214071 106934
rect 252277 106931 252343 106934
rect 177246 106796 177252 106860
rect 177316 106858 177322 106860
rect 195421 106858 195487 106861
rect 177316 106856 195487 106858
rect 177316 106800 195426 106856
rect 195482 106800 195487 106856
rect 306741 106858 306807 106861
rect 306741 106856 310040 106858
rect 177316 106798 195487 106800
rect 177316 106796 177322 106798
rect 195421 106795 195487 106798
rect 213913 106450 213979 106453
rect 217182 106450 217242 106828
rect 306741 106800 306746 106856
rect 306802 106800 310040 106856
rect 306741 106798 310040 106800
rect 306741 106795 306807 106798
rect 252369 106586 252435 106589
rect 248952 106584 252435 106586
rect 248952 106528 252374 106584
rect 252430 106528 252435 106584
rect 248952 106526 252435 106528
rect 252369 106523 252435 106526
rect 213913 106448 217242 106450
rect 213913 106392 213918 106448
rect 213974 106392 217242 106448
rect 213913 106390 217242 106392
rect 305913 106450 305979 106453
rect 305913 106448 310040 106450
rect 305913 106392 305918 106448
rect 305974 106392 310040 106448
rect 305913 106390 310040 106392
rect 213913 106387 213979 106390
rect 305913 106387 305979 106390
rect 328494 106314 328500 106316
rect 321908 106254 328500 106314
rect 328494 106252 328500 106254
rect 328564 106252 328570 106316
rect 213913 105770 213979 105773
rect 217182 105770 217242 106148
rect 251173 106042 251239 106045
rect 248952 106040 251239 106042
rect 248952 105984 251178 106040
rect 251234 105984 251239 106040
rect 248952 105982 251239 105984
rect 251173 105979 251239 105982
rect 307569 105906 307635 105909
rect 307569 105904 310040 105906
rect 307569 105848 307574 105904
rect 307630 105848 310040 105904
rect 307569 105846 310040 105848
rect 307569 105843 307635 105846
rect 213913 105768 217242 105770
rect 213913 105712 213918 105768
rect 213974 105712 217242 105768
rect 213913 105710 217242 105712
rect 213913 105707 213979 105710
rect 252461 105634 252527 105637
rect 248952 105632 252527 105634
rect 173014 105164 173020 105228
rect 173084 105226 173090 105228
rect 217182 105226 217242 105604
rect 248952 105576 252466 105632
rect 252522 105576 252527 105632
rect 248952 105574 252527 105576
rect 252461 105571 252527 105574
rect 324313 105498 324379 105501
rect 321908 105496 324379 105498
rect 309550 105394 310132 105454
rect 321908 105440 324318 105496
rect 324374 105440 324379 105496
rect 321908 105438 324379 105440
rect 324313 105435 324379 105438
rect 305637 105362 305703 105365
rect 309550 105362 309610 105394
rect 305637 105360 309610 105362
rect 305637 105304 305642 105360
rect 305698 105304 309610 105360
rect 305637 105302 309610 105304
rect 305637 105299 305703 105302
rect 173084 105166 217242 105226
rect 173084 105164 173090 105166
rect 214598 105028 214604 105092
rect 214668 105090 214674 105092
rect 252185 105090 252251 105093
rect 214668 105030 217242 105090
rect 248952 105088 252251 105090
rect 248952 105032 252190 105088
rect 252246 105032 252251 105088
rect 248952 105030 252251 105032
rect 214668 105028 214674 105030
rect 217182 104924 217242 105030
rect 252185 105027 252251 105030
rect 307661 105090 307727 105093
rect 307661 105088 310040 105090
rect 307661 105032 307666 105088
rect 307722 105032 310040 105088
rect 307661 105030 310040 105032
rect 307661 105027 307727 105030
rect 324313 104818 324379 104821
rect 321908 104816 324379 104818
rect 321908 104760 324318 104816
rect 324374 104760 324379 104816
rect 321908 104758 324379 104760
rect 324313 104755 324379 104758
rect 251766 104682 251772 104684
rect 248952 104622 251772 104682
rect 251766 104620 251772 104622
rect 251836 104620 251842 104684
rect 307477 104682 307543 104685
rect 307477 104680 310040 104682
rect 307477 104624 307482 104680
rect 307538 104624 310040 104680
rect 307477 104622 310040 104624
rect 307477 104619 307543 104622
rect 307569 104274 307635 104277
rect 307569 104272 310040 104274
rect 214005 104002 214071 104005
rect 217182 104002 217242 104244
rect 307569 104216 307574 104272
rect 307630 104216 310040 104272
rect 307569 104214 310040 104216
rect 307569 104211 307635 104214
rect 252461 104138 252527 104141
rect 248952 104136 252527 104138
rect 248952 104080 252466 104136
rect 252522 104080 252527 104136
rect 248952 104078 252527 104080
rect 252461 104075 252527 104078
rect 325601 104002 325667 104005
rect 214005 104000 217242 104002
rect 214005 103944 214010 104000
rect 214066 103944 217242 104000
rect 214005 103942 217242 103944
rect 321908 104000 325667 104002
rect 321908 103944 325606 104000
rect 325662 103944 325667 104000
rect 321908 103942 325667 103944
rect 214005 103939 214071 103942
rect 325601 103939 325667 103942
rect 307661 103866 307727 103869
rect 307661 103864 310040 103866
rect 307661 103808 307666 103864
rect 307722 103808 310040 103864
rect 307661 103806 310040 103808
rect 307661 103803 307727 103806
rect 213913 103730 213979 103733
rect 252093 103730 252159 103733
rect 213913 103728 217242 103730
rect 213913 103672 213918 103728
rect 213974 103672 217242 103728
rect 213913 103670 217242 103672
rect 248952 103728 252159 103730
rect 248952 103672 252098 103728
rect 252154 103672 252159 103728
rect 248952 103670 252159 103672
rect 213913 103667 213979 103670
rect 217182 103564 217242 103670
rect 252093 103667 252159 103670
rect 307477 103458 307543 103461
rect 307477 103456 310040 103458
rect 307477 103400 307482 103456
rect 307538 103400 310040 103456
rect 307477 103398 310040 103400
rect 307477 103395 307543 103398
rect 252461 103186 252527 103189
rect 324313 103186 324379 103189
rect 248952 103184 252527 103186
rect 248952 103128 252466 103184
rect 252522 103128 252527 103184
rect 248952 103126 252527 103128
rect 321908 103184 324379 103186
rect 321908 103128 324318 103184
rect 324374 103128 324379 103184
rect 321908 103126 324379 103128
rect 252461 103123 252527 103126
rect 324313 103123 324379 103126
rect 307569 103050 307635 103053
rect 307569 103048 310040 103050
rect 307569 102992 307574 103048
rect 307630 102992 310040 103048
rect 307569 102990 310040 102992
rect 307569 102987 307635 102990
rect 214005 102506 214071 102509
rect 217182 102506 217242 102884
rect 252185 102778 252251 102781
rect 248952 102776 252251 102778
rect 248952 102720 252190 102776
rect 252246 102720 252251 102776
rect 248952 102718 252251 102720
rect 252185 102715 252251 102718
rect 214005 102504 217242 102506
rect 214005 102448 214010 102504
rect 214066 102448 217242 102504
rect 214005 102446 217242 102448
rect 307661 102506 307727 102509
rect 324497 102506 324563 102509
rect 307661 102504 310040 102506
rect 307661 102448 307666 102504
rect 307722 102448 310040 102504
rect 307661 102446 310040 102448
rect 321908 102504 324563 102506
rect 321908 102448 324502 102504
rect 324558 102448 324563 102504
rect 321908 102446 324563 102448
rect 214005 102443 214071 102446
rect 307661 102443 307727 102446
rect 324497 102443 324563 102446
rect 66069 102370 66135 102373
rect 68142 102370 68816 102376
rect 66069 102368 68816 102370
rect 66069 102312 66074 102368
rect 66130 102316 68816 102368
rect 213913 102370 213979 102373
rect 213913 102368 217242 102370
rect 66130 102312 68202 102316
rect 66069 102310 68202 102312
rect 213913 102312 213918 102368
rect 213974 102312 217242 102368
rect 213913 102310 217242 102312
rect 66069 102307 66135 102310
rect 213913 102307 213979 102310
rect 217182 102204 217242 102310
rect 252369 102234 252435 102237
rect 248952 102232 252435 102234
rect 248952 102176 252374 102232
rect 252430 102176 252435 102232
rect 248952 102174 252435 102176
rect 252369 102171 252435 102174
rect 307569 102098 307635 102101
rect 307569 102096 310040 102098
rect 307569 102040 307574 102096
rect 307630 102040 310040 102096
rect 307569 102038 310040 102040
rect 307569 102035 307635 102038
rect 254526 101826 254532 101828
rect 248952 101766 254532 101826
rect 254526 101764 254532 101766
rect 254596 101764 254602 101828
rect 309550 101586 310132 101646
rect 214005 101282 214071 101285
rect 217182 101282 217242 101524
rect 252277 101418 252343 101421
rect 248952 101416 252343 101418
rect 248952 101360 252282 101416
rect 252338 101360 252343 101416
rect 248952 101358 252343 101360
rect 252277 101355 252343 101358
rect 214005 101280 217242 101282
rect 214005 101224 214010 101280
rect 214066 101224 217242 101280
rect 214005 101222 217242 101224
rect 214005 101219 214071 101222
rect 213913 101146 213979 101149
rect 305729 101146 305795 101149
rect 309550 101146 309610 101586
rect 213913 101144 217242 101146
rect 213913 101088 213918 101144
rect 213974 101088 217242 101144
rect 213913 101086 217242 101088
rect 213913 101083 213979 101086
rect 217182 100980 217242 101086
rect 305729 101144 309610 101146
rect 305729 101088 305734 101144
rect 305790 101088 309610 101144
rect 305729 101086 309610 101088
rect 309734 101178 310132 101238
rect 305729 101083 305795 101086
rect 307477 101010 307543 101013
rect 309734 101010 309794 101178
rect 307477 101008 309794 101010
rect 307477 100952 307482 101008
rect 307538 100952 309794 101008
rect 307477 100950 309794 100952
rect 321878 101010 321938 101660
rect 338246 101010 338252 101012
rect 321878 100950 338252 101010
rect 307477 100947 307543 100950
rect 338246 100948 338252 100950
rect 338316 100948 338322 101012
rect 252461 100874 252527 100877
rect 248952 100872 252527 100874
rect 248952 100816 252466 100872
rect 252522 100816 252527 100872
rect 248952 100814 252527 100816
rect 252461 100811 252527 100814
rect 307661 100874 307727 100877
rect 307661 100872 310040 100874
rect 307661 100816 307666 100872
rect 307722 100816 310040 100872
rect 307661 100814 310040 100816
rect 307661 100811 307727 100814
rect 67633 100738 67699 100741
rect 68142 100738 68816 100744
rect 67633 100736 68816 100738
rect 67633 100680 67638 100736
rect 67694 100684 68816 100736
rect 67694 100680 68202 100684
rect 67633 100678 68202 100680
rect 67633 100675 67699 100678
rect 321326 100469 321386 100844
rect 252461 100466 252527 100469
rect 248952 100464 252527 100466
rect 248952 100408 252466 100464
rect 252522 100408 252527 100464
rect 248952 100406 252527 100408
rect 252461 100403 252527 100406
rect 307569 100466 307635 100469
rect 307569 100464 310040 100466
rect 307569 100408 307574 100464
rect 307630 100408 310040 100464
rect 307569 100406 310040 100408
rect 321277 100464 321386 100469
rect 321277 100408 321282 100464
rect 321338 100408 321386 100464
rect 321277 100406 321386 100408
rect 307569 100403 307635 100406
rect 321277 100403 321343 100406
rect 214097 99786 214163 99789
rect 217182 99786 217242 100300
rect 324313 100194 324379 100197
rect 321908 100192 324379 100194
rect 321908 100136 324318 100192
rect 324374 100136 324379 100192
rect 321908 100134 324379 100136
rect 324313 100131 324379 100134
rect 306741 100058 306807 100061
rect 306741 100056 310040 100058
rect 306741 100000 306746 100056
rect 306802 100000 310040 100056
rect 306741 99998 310040 100000
rect 306741 99995 306807 99998
rect 252369 99922 252435 99925
rect 248952 99920 252435 99922
rect 248952 99864 252374 99920
rect 252430 99864 252435 99920
rect 248952 99862 252435 99864
rect 252369 99859 252435 99862
rect 214097 99784 217242 99786
rect 214097 99728 214102 99784
rect 214158 99728 217242 99784
rect 214097 99726 217242 99728
rect 214097 99723 214163 99726
rect 307661 99650 307727 99653
rect 307661 99648 310040 99650
rect 170254 99452 170260 99516
rect 170324 99514 170330 99516
rect 170324 99454 216874 99514
rect 170324 99452 170330 99454
rect 216814 99378 216874 99454
rect 217366 99378 217426 99620
rect 307661 99592 307666 99648
rect 307722 99592 310040 99648
rect 307661 99590 310040 99592
rect 307661 99587 307727 99590
rect 252277 99514 252343 99517
rect 248952 99512 252343 99514
rect 248952 99456 252282 99512
rect 252338 99456 252343 99512
rect 248952 99454 252343 99456
rect 252277 99451 252343 99454
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 216814 99318 217426 99378
rect 583520 99364 584960 99454
rect 307569 99106 307635 99109
rect 307569 99104 310040 99106
rect 307569 99048 307574 99104
rect 307630 99048 310040 99104
rect 307569 99046 310040 99048
rect 307569 99043 307635 99046
rect 253197 98970 253263 98973
rect 248952 98968 253263 98970
rect 214005 98426 214071 98429
rect 217182 98426 217242 98940
rect 248952 98912 253202 98968
rect 253258 98912 253263 98968
rect 248952 98910 253263 98912
rect 253197 98907 253263 98910
rect 321369 98834 321435 98837
rect 321510 98834 321570 99348
rect 321369 98832 321570 98834
rect 321369 98776 321374 98832
rect 321430 98776 321570 98832
rect 321369 98774 321570 98776
rect 321369 98771 321435 98774
rect 307109 98698 307175 98701
rect 307109 98696 310040 98698
rect 307109 98640 307114 98696
rect 307170 98640 310040 98696
rect 307109 98638 310040 98640
rect 307109 98635 307175 98638
rect 252461 98562 252527 98565
rect 324589 98562 324655 98565
rect 248952 98560 252527 98562
rect 248952 98504 252466 98560
rect 252522 98504 252527 98560
rect 248952 98502 252527 98504
rect 321908 98560 324655 98562
rect 321908 98504 324594 98560
rect 324650 98504 324655 98560
rect 321908 98502 324655 98504
rect 252461 98499 252527 98502
rect 324589 98499 324655 98502
rect 214005 98424 217242 98426
rect 214005 98368 214010 98424
rect 214066 98368 217242 98424
rect 214005 98366 217242 98368
rect 214005 98363 214071 98366
rect 307661 98290 307727 98293
rect 307661 98288 310040 98290
rect 213913 98018 213979 98021
rect 217366 98018 217426 98260
rect 307661 98232 307666 98288
rect 307722 98232 310040 98288
rect 307661 98230 310040 98232
rect 307661 98227 307727 98230
rect 252369 98018 252435 98021
rect 213913 98016 217426 98018
rect 213913 97960 213918 98016
rect 213974 97960 217426 98016
rect 213913 97958 217426 97960
rect 248952 98016 252435 98018
rect 248952 97960 252374 98016
rect 252430 97960 252435 98016
rect 248952 97958 252435 97960
rect 213913 97955 213979 97958
rect 252369 97955 252435 97958
rect 307661 97882 307727 97885
rect 307661 97880 310040 97882
rect 307661 97824 307666 97880
rect 307722 97824 310040 97880
rect 307661 97822 310040 97824
rect 307661 97819 307727 97822
rect -960 97610 480 97700
rect 3509 97610 3575 97613
rect 252185 97610 252251 97613
rect -960 97608 3575 97610
rect -960 97552 3514 97608
rect 3570 97552 3575 97608
rect 248952 97608 252251 97610
rect -960 97550 3575 97552
rect -960 97460 480 97550
rect 3509 97547 3575 97550
rect 214414 97004 214420 97068
rect 214484 97066 214490 97068
rect 217182 97066 217242 97580
rect 248952 97552 252190 97608
rect 252246 97552 252251 97608
rect 248952 97550 252251 97552
rect 252185 97547 252251 97550
rect 306925 97474 306991 97477
rect 306925 97472 310040 97474
rect 306925 97416 306930 97472
rect 306986 97416 310040 97472
rect 306925 97414 310040 97416
rect 306925 97411 306991 97414
rect 321510 97341 321570 97852
rect 321510 97336 321619 97341
rect 321510 97280 321558 97336
rect 321614 97280 321619 97336
rect 321510 97278 321619 97280
rect 321553 97275 321619 97278
rect 251265 97066 251331 97069
rect 252461 97066 252527 97069
rect 214484 97006 217242 97066
rect 248952 97064 252527 97066
rect 248952 97008 251270 97064
rect 251326 97008 252466 97064
rect 252522 97008 252527 97064
rect 248952 97006 252527 97008
rect 214484 97004 214490 97006
rect 251265 97003 251331 97006
rect 252461 97003 252527 97006
rect 307150 97004 307156 97068
rect 307220 97066 307226 97068
rect 324446 97066 324452 97068
rect 307220 97006 310040 97066
rect 321908 97006 324452 97066
rect 307220 97004 307226 97006
rect 324446 97004 324452 97006
rect 324516 97004 324522 97068
rect 214557 96658 214623 96661
rect 217182 96658 217242 96900
rect 249149 96658 249215 96661
rect 262070 96658 262076 96660
rect 214557 96656 217242 96658
rect 214557 96600 214562 96656
rect 214618 96600 217242 96656
rect 214557 96598 217242 96600
rect 248952 96656 262076 96658
rect 248952 96600 249154 96656
rect 249210 96600 262076 96656
rect 248952 96598 262076 96600
rect 214557 96595 214623 96598
rect 249149 96595 249215 96598
rect 262070 96596 262076 96598
rect 262140 96596 262146 96660
rect 307661 96658 307727 96661
rect 321461 96658 321527 96661
rect 307661 96656 310040 96658
rect 307661 96600 307666 96656
rect 307722 96600 310040 96656
rect 307661 96598 310040 96600
rect 321461 96656 321570 96658
rect 321461 96600 321466 96656
rect 321522 96600 321570 96656
rect 307661 96595 307727 96598
rect 321461 96595 321570 96600
rect 321510 96356 321570 96595
rect 214741 95842 214807 95845
rect 217182 95842 217242 96356
rect 251173 96250 251239 96253
rect 248860 96248 251239 96250
rect 248860 96192 251178 96248
rect 251234 96192 251239 96248
rect 248860 96190 251239 96192
rect 251173 96187 251239 96190
rect 306925 96250 306991 96253
rect 306925 96248 310132 96250
rect 306925 96192 306930 96248
rect 306986 96192 310132 96248
rect 306925 96190 310132 96192
rect 306925 96187 306991 96190
rect 214741 95840 217242 95842
rect 214741 95784 214746 95840
rect 214802 95784 217242 95840
rect 214741 95782 217242 95784
rect 214741 95779 214807 95782
rect 178677 95162 178743 95165
rect 321369 95162 321435 95165
rect 178677 95160 321435 95162
rect 178677 95104 178682 95160
rect 178738 95104 321374 95160
rect 321430 95104 321435 95160
rect 178677 95102 321435 95104
rect 178677 95099 178743 95102
rect 321369 95099 321435 95102
rect 66161 94890 66227 94893
rect 173014 94890 173020 94892
rect 66161 94888 173020 94890
rect 66161 94832 66166 94888
rect 66222 94832 173020 94888
rect 66161 94830 173020 94832
rect 66161 94827 66227 94830
rect 173014 94828 173020 94830
rect 173084 94828 173090 94892
rect 129365 94756 129431 94757
rect 106222 94692 106228 94756
rect 106292 94754 106298 94756
rect 106608 94754 106614 94756
rect 106292 94694 106614 94754
rect 106292 94692 106298 94694
rect 106608 94692 106614 94694
rect 106678 94692 106684 94756
rect 129320 94692 129326 94756
rect 129390 94754 129431 94756
rect 151721 94756 151787 94757
rect 151721 94754 151766 94756
rect 129390 94752 129482 94754
rect 129426 94696 129482 94752
rect 129390 94694 129482 94696
rect 151674 94752 151766 94754
rect 151674 94696 151726 94752
rect 151674 94694 151766 94696
rect 129390 94692 129431 94694
rect 129365 94691 129431 94692
rect 151721 94692 151766 94694
rect 151830 94692 151836 94756
rect 151721 94691 151787 94692
rect 111926 93876 111932 93940
rect 111996 93938 112002 93940
rect 169150 93938 169156 93940
rect 111996 93878 169156 93938
rect 111996 93876 112002 93878
rect 169150 93876 169156 93878
rect 169220 93876 169226 93940
rect 67449 93802 67515 93805
rect 214598 93802 214604 93804
rect 67449 93800 214604 93802
rect 67449 93744 67454 93800
rect 67510 93744 214604 93800
rect 67449 93742 214604 93744
rect 67449 93739 67515 93742
rect 214598 93740 214604 93742
rect 214668 93740 214674 93804
rect 85665 93668 85731 93669
rect 115473 93668 115539 93669
rect 120625 93668 120691 93669
rect 135713 93668 135779 93669
rect 151721 93668 151787 93669
rect 85614 93666 85620 93668
rect 85574 93606 85620 93666
rect 85684 93664 85731 93668
rect 115422 93666 115428 93668
rect 85726 93608 85731 93664
rect 85614 93604 85620 93606
rect 85684 93604 85731 93608
rect 115382 93606 115428 93666
rect 115492 93664 115539 93668
rect 120574 93666 120580 93668
rect 115534 93608 115539 93664
rect 115422 93604 115428 93606
rect 115492 93604 115539 93608
rect 120534 93606 120580 93666
rect 120644 93664 120691 93668
rect 135662 93666 135668 93668
rect 120686 93608 120691 93664
rect 120574 93604 120580 93606
rect 120644 93604 120691 93608
rect 135622 93606 135668 93666
rect 135732 93664 135779 93668
rect 135774 93608 135779 93664
rect 135662 93604 135668 93606
rect 135732 93604 135779 93608
rect 151670 93604 151676 93668
rect 151740 93666 151787 93668
rect 195329 93666 195395 93669
rect 324446 93666 324452 93668
rect 151740 93664 151832 93666
rect 151782 93608 151832 93664
rect 151740 93606 151832 93608
rect 195329 93664 324452 93666
rect 195329 93608 195334 93664
rect 195390 93608 324452 93664
rect 195329 93606 324452 93608
rect 151740 93604 151787 93606
rect 85665 93603 85731 93604
rect 115473 93603 115539 93604
rect 120625 93603 120691 93604
rect 135713 93603 135779 93604
rect 151721 93603 151787 93604
rect 195329 93603 195395 93606
rect 324446 93604 324452 93606
rect 324516 93604 324522 93668
rect 61929 93530 61995 93533
rect 199561 93530 199627 93533
rect 61929 93528 199627 93530
rect 61929 93472 61934 93528
rect 61990 93472 199566 93528
rect 199622 93472 199627 93528
rect 61929 93470 199627 93472
rect 61929 93467 61995 93470
rect 199561 93467 199627 93470
rect 103278 93196 103284 93260
rect 103348 93258 103354 93260
rect 103421 93258 103487 93261
rect 110321 93260 110387 93261
rect 113817 93260 113883 93261
rect 128169 93260 128235 93261
rect 110270 93258 110276 93260
rect 103348 93256 103487 93258
rect 103348 93200 103426 93256
rect 103482 93200 103487 93256
rect 103348 93198 103487 93200
rect 110230 93198 110276 93258
rect 110340 93256 110387 93260
rect 113766 93258 113772 93260
rect 110382 93200 110387 93256
rect 103348 93196 103354 93198
rect 103421 93195 103487 93198
rect 110270 93196 110276 93198
rect 110340 93196 110387 93200
rect 113726 93198 113772 93258
rect 113836 93256 113883 93260
rect 128118 93258 128124 93260
rect 113878 93200 113883 93256
rect 113766 93196 113772 93198
rect 113836 93196 113883 93200
rect 128078 93198 128124 93258
rect 128188 93256 128235 93260
rect 128230 93200 128235 93256
rect 128118 93196 128124 93198
rect 128188 93196 128235 93200
rect 110321 93195 110387 93196
rect 113817 93195 113883 93196
rect 128169 93195 128235 93196
rect 74809 92444 74875 92445
rect 88977 92444 89043 92445
rect 95049 92444 95115 92445
rect 74758 92442 74764 92444
rect 74718 92382 74764 92442
rect 74828 92440 74875 92444
rect 88926 92442 88932 92444
rect 74870 92384 74875 92440
rect 74758 92380 74764 92382
rect 74828 92380 74875 92384
rect 88886 92382 88932 92442
rect 88996 92440 89043 92444
rect 94998 92442 95004 92444
rect 89038 92384 89043 92440
rect 88926 92380 88932 92382
rect 88996 92380 89043 92384
rect 94958 92382 95004 92442
rect 95068 92440 95115 92444
rect 95110 92384 95115 92440
rect 94998 92380 95004 92382
rect 95068 92380 95115 92384
rect 101806 92380 101812 92444
rect 101876 92442 101882 92444
rect 102041 92442 102107 92445
rect 105537 92444 105603 92445
rect 105486 92442 105492 92444
rect 101876 92440 102107 92442
rect 101876 92384 102046 92440
rect 102102 92384 102107 92440
rect 101876 92382 102107 92384
rect 105446 92382 105492 92442
rect 105556 92440 105603 92444
rect 105598 92384 105603 92440
rect 101876 92380 101882 92382
rect 74809 92379 74875 92380
rect 88977 92379 89043 92380
rect 95049 92379 95115 92380
rect 102041 92379 102107 92382
rect 105486 92380 105492 92382
rect 105556 92380 105603 92384
rect 106222 92380 106228 92444
rect 106292 92442 106298 92444
rect 106641 92442 106707 92445
rect 116761 92444 116827 92445
rect 116710 92442 116716 92444
rect 106292 92440 106707 92442
rect 106292 92384 106646 92440
rect 106702 92384 106707 92440
rect 106292 92382 106707 92384
rect 116670 92382 116716 92442
rect 116780 92440 116827 92444
rect 116822 92384 116827 92440
rect 106292 92380 106298 92382
rect 105537 92379 105603 92380
rect 106641 92379 106707 92382
rect 116710 92380 116716 92382
rect 116780 92380 116827 92384
rect 116761 92379 116827 92380
rect 124029 92444 124095 92445
rect 124029 92440 124076 92444
rect 124140 92442 124146 92444
rect 124029 92384 124034 92440
rect 124029 92380 124076 92384
rect 124140 92382 124186 92442
rect 124140 92380 124146 92382
rect 125726 92380 125732 92444
rect 125796 92442 125802 92444
rect 126697 92442 126763 92445
rect 134425 92444 134491 92445
rect 134374 92442 134380 92444
rect 125796 92440 126763 92442
rect 125796 92384 126702 92440
rect 126758 92384 126763 92440
rect 125796 92382 126763 92384
rect 134334 92382 134380 92442
rect 134444 92440 134491 92444
rect 134486 92384 134491 92440
rect 125796 92380 125802 92382
rect 124029 92379 124095 92380
rect 126697 92379 126763 92382
rect 134374 92380 134380 92382
rect 134444 92380 134491 92384
rect 152038 92380 152044 92444
rect 152108 92442 152114 92444
rect 153009 92442 153075 92445
rect 152108 92440 153075 92442
rect 152108 92384 153014 92440
rect 153070 92384 153075 92440
rect 152108 92382 153075 92384
rect 152108 92380 152114 92382
rect 134425 92379 134491 92380
rect 153009 92379 153075 92382
rect 114318 92244 114324 92308
rect 114388 92306 114394 92308
rect 178953 92306 179019 92309
rect 114388 92304 179019 92306
rect 114388 92248 178958 92304
rect 179014 92248 179019 92304
rect 114388 92246 179019 92248
rect 114388 92244 114394 92246
rect 178953 92243 179019 92246
rect 126697 92036 126763 92037
rect 126646 92034 126652 92036
rect 126606 91974 126652 92034
rect 126716 92032 126763 92036
rect 126758 91976 126763 92032
rect 126646 91972 126652 91974
rect 126716 91972 126763 91976
rect 126697 91971 126763 91972
rect 105670 91700 105676 91764
rect 105740 91762 105746 91764
rect 106089 91762 106155 91765
rect 105740 91760 106155 91762
rect 105740 91704 106094 91760
rect 106150 91704 106155 91760
rect 105740 91702 106155 91704
rect 105740 91700 105746 91702
rect 106089 91699 106155 91702
rect 114870 91700 114876 91764
rect 114940 91762 114946 91764
rect 115565 91762 115631 91765
rect 114940 91760 115631 91762
rect 114940 91704 115570 91760
rect 115626 91704 115631 91760
rect 114940 91702 115631 91704
rect 114940 91700 114946 91702
rect 115565 91699 115631 91702
rect 124438 91564 124444 91628
rect 124508 91626 124514 91628
rect 125409 91626 125475 91629
rect 124508 91624 125475 91626
rect 124508 91568 125414 91624
rect 125470 91568 125475 91624
rect 124508 91566 125475 91568
rect 124508 91564 124514 91566
rect 125409 91563 125475 91566
rect 126462 91564 126468 91628
rect 126532 91626 126538 91628
rect 126881 91626 126947 91629
rect 126532 91624 126947 91626
rect 126532 91568 126886 91624
rect 126942 91568 126947 91624
rect 126532 91566 126947 91568
rect 126532 91564 126538 91566
rect 126881 91563 126947 91566
rect 122833 91492 122899 91493
rect 122782 91428 122788 91492
rect 122852 91490 122899 91492
rect 122852 91488 122944 91490
rect 122894 91432 122944 91488
rect 122852 91430 122944 91432
rect 122852 91428 122899 91430
rect 122833 91427 122899 91428
rect 98494 91292 98500 91356
rect 98564 91354 98570 91356
rect 99189 91354 99255 91357
rect 98564 91352 99255 91354
rect 98564 91296 99194 91352
rect 99250 91296 99255 91352
rect 98564 91294 99255 91296
rect 98564 91292 98570 91294
rect 99189 91291 99255 91294
rect 100886 91292 100892 91356
rect 100956 91354 100962 91356
rect 101857 91354 101923 91357
rect 100956 91352 101923 91354
rect 100956 91296 101862 91352
rect 101918 91296 101923 91352
rect 100956 91294 101923 91296
rect 100956 91292 100962 91294
rect 101857 91291 101923 91294
rect 104198 91292 104204 91356
rect 104268 91354 104274 91356
rect 104801 91354 104867 91357
rect 104268 91352 104867 91354
rect 104268 91296 104806 91352
rect 104862 91296 104867 91352
rect 104268 91294 104867 91296
rect 104268 91292 104274 91294
rect 104801 91291 104867 91294
rect 108062 91292 108068 91356
rect 108132 91354 108138 91356
rect 108205 91354 108271 91357
rect 109585 91356 109651 91357
rect 118233 91356 118299 91357
rect 109534 91354 109540 91356
rect 108132 91352 108271 91354
rect 108132 91296 108210 91352
rect 108266 91296 108271 91352
rect 108132 91294 108271 91296
rect 109494 91294 109540 91354
rect 109604 91352 109651 91356
rect 118182 91354 118188 91356
rect 109646 91296 109651 91352
rect 108132 91292 108138 91294
rect 108205 91291 108271 91294
rect 109534 91292 109540 91294
rect 109604 91292 109651 91296
rect 118142 91294 118188 91354
rect 118252 91352 118299 91356
rect 118294 91296 118299 91352
rect 118182 91292 118188 91294
rect 118252 91292 118299 91296
rect 119286 91292 119292 91356
rect 119356 91354 119362 91356
rect 119889 91354 119955 91357
rect 119356 91352 119955 91354
rect 119356 91296 119894 91352
rect 119950 91296 119955 91352
rect 119356 91294 119955 91296
rect 119356 91292 119362 91294
rect 109585 91291 109651 91292
rect 118233 91291 118299 91292
rect 119889 91291 119955 91294
rect 121678 91292 121684 91356
rect 121748 91354 121754 91356
rect 122649 91354 122715 91357
rect 121748 91352 122715 91354
rect 121748 91296 122654 91352
rect 122710 91296 122715 91352
rect 121748 91294 122715 91296
rect 121748 91292 121754 91294
rect 122649 91291 122715 91294
rect 84326 91156 84332 91220
rect 84396 91218 84402 91220
rect 85481 91218 85547 91221
rect 84396 91216 85547 91218
rect 84396 91160 85486 91216
rect 85542 91160 85547 91216
rect 84396 91158 85547 91160
rect 84396 91156 84402 91158
rect 85481 91155 85547 91158
rect 86718 91156 86724 91220
rect 86788 91218 86794 91220
rect 86861 91218 86927 91221
rect 88057 91220 88123 91221
rect 88006 91218 88012 91220
rect 86788 91216 86927 91218
rect 86788 91160 86866 91216
rect 86922 91160 86927 91216
rect 86788 91158 86927 91160
rect 87966 91158 88012 91218
rect 88076 91216 88123 91220
rect 88118 91160 88123 91216
rect 86788 91156 86794 91158
rect 86861 91155 86927 91158
rect 88006 91156 88012 91158
rect 88076 91156 88123 91160
rect 90214 91156 90220 91220
rect 90284 91218 90290 91220
rect 90725 91218 90791 91221
rect 90284 91216 90791 91218
rect 90284 91160 90730 91216
rect 90786 91160 90791 91216
rect 90284 91158 90791 91160
rect 90284 91156 90290 91158
rect 88057 91155 88123 91156
rect 90725 91155 90791 91158
rect 91318 91156 91324 91220
rect 91388 91218 91394 91220
rect 92381 91218 92447 91221
rect 91388 91216 92447 91218
rect 91388 91160 92386 91216
rect 92442 91160 92447 91216
rect 91388 91158 92447 91160
rect 91388 91156 91394 91158
rect 92381 91155 92447 91158
rect 92606 91156 92612 91220
rect 92676 91218 92682 91220
rect 93761 91218 93827 91221
rect 92676 91216 93827 91218
rect 92676 91160 93766 91216
rect 93822 91160 93827 91216
rect 92676 91158 93827 91160
rect 92676 91156 92682 91158
rect 93761 91155 93827 91158
rect 93894 91156 93900 91220
rect 93964 91218 93970 91220
rect 95141 91218 95207 91221
rect 93964 91216 95207 91218
rect 93964 91160 95146 91216
rect 95202 91160 95207 91216
rect 93964 91158 95207 91160
rect 93964 91156 93970 91158
rect 95141 91155 95207 91158
rect 96286 91156 96292 91220
rect 96356 91218 96362 91220
rect 96521 91218 96587 91221
rect 96356 91216 96587 91218
rect 96356 91160 96526 91216
rect 96582 91160 96587 91216
rect 96356 91158 96587 91160
rect 96356 91156 96362 91158
rect 96521 91155 96587 91158
rect 96654 91156 96660 91220
rect 96724 91218 96730 91220
rect 97073 91218 97139 91221
rect 96724 91216 97139 91218
rect 96724 91160 97078 91216
rect 97134 91160 97139 91216
rect 96724 91158 97139 91160
rect 96724 91156 96730 91158
rect 97073 91155 97139 91158
rect 97206 91156 97212 91220
rect 97276 91218 97282 91220
rect 97901 91218 97967 91221
rect 97276 91216 97967 91218
rect 97276 91160 97906 91216
rect 97962 91160 97967 91216
rect 97276 91158 97967 91160
rect 97276 91156 97282 91158
rect 97901 91155 97967 91158
rect 98126 91156 98132 91220
rect 98196 91156 98202 91220
rect 99046 91156 99052 91220
rect 99116 91218 99122 91220
rect 99281 91218 99347 91221
rect 99116 91216 99347 91218
rect 99116 91160 99286 91216
rect 99342 91160 99347 91216
rect 99116 91158 99347 91160
rect 99116 91156 99122 91158
rect 98134 91082 98194 91156
rect 99281 91155 99347 91158
rect 99966 91156 99972 91220
rect 100036 91218 100042 91220
rect 100201 91218 100267 91221
rect 100036 91216 100267 91218
rect 100036 91160 100206 91216
rect 100262 91160 100267 91216
rect 100036 91158 100267 91160
rect 100036 91156 100042 91158
rect 100201 91155 100267 91158
rect 100518 91156 100524 91220
rect 100588 91218 100594 91220
rect 100661 91218 100727 91221
rect 101949 91220 102015 91221
rect 101949 91218 101996 91220
rect 100588 91216 100727 91218
rect 100588 91160 100666 91216
rect 100722 91160 100727 91216
rect 100588 91158 100727 91160
rect 101904 91216 101996 91218
rect 101904 91160 101954 91216
rect 101904 91158 101996 91160
rect 100588 91156 100594 91158
rect 100661 91155 100727 91158
rect 101949 91156 101996 91158
rect 102060 91156 102066 91220
rect 102726 91156 102732 91220
rect 102796 91218 102802 91220
rect 102961 91218 103027 91221
rect 102796 91216 103027 91218
rect 102796 91160 102966 91216
rect 103022 91160 103027 91216
rect 102796 91158 103027 91160
rect 102796 91156 102802 91158
rect 101949 91155 102015 91156
rect 102961 91155 103027 91158
rect 104566 91156 104572 91220
rect 104636 91218 104642 91220
rect 104709 91218 104775 91221
rect 104636 91216 104775 91218
rect 104636 91160 104714 91216
rect 104770 91160 104775 91216
rect 104636 91158 104775 91160
rect 104636 91156 104642 91158
rect 104709 91155 104775 91158
rect 106590 91156 106596 91220
rect 106660 91218 106666 91220
rect 107193 91218 107259 91221
rect 106660 91216 107259 91218
rect 106660 91160 107198 91216
rect 107254 91160 107259 91216
rect 106660 91158 107259 91160
rect 106660 91156 106666 91158
rect 107193 91155 107259 91158
rect 107694 91156 107700 91220
rect 107764 91218 107770 91220
rect 108481 91218 108547 91221
rect 107764 91216 108547 91218
rect 107764 91160 108486 91216
rect 108542 91160 108547 91216
rect 107764 91158 108547 91160
rect 107764 91156 107770 91158
rect 108481 91155 108547 91158
rect 109166 91156 109172 91220
rect 109236 91218 109242 91220
rect 110137 91218 110203 91221
rect 110689 91220 110755 91221
rect 110638 91218 110644 91220
rect 109236 91216 110203 91218
rect 109236 91160 110142 91216
rect 110198 91160 110203 91216
rect 109236 91158 110203 91160
rect 110598 91158 110644 91218
rect 110708 91216 110755 91220
rect 110750 91160 110755 91216
rect 109236 91156 109242 91158
rect 110137 91155 110203 91158
rect 110638 91156 110644 91158
rect 110708 91156 110755 91160
rect 111190 91156 111196 91220
rect 111260 91218 111266 91220
rect 111701 91218 111767 91221
rect 111260 91216 111767 91218
rect 111260 91160 111706 91216
rect 111762 91160 111767 91216
rect 111260 91158 111767 91160
rect 111260 91156 111266 91158
rect 110689 91155 110755 91156
rect 111701 91155 111767 91158
rect 112294 91156 112300 91220
rect 112364 91218 112370 91220
rect 112529 91218 112595 91221
rect 112364 91216 112595 91218
rect 112364 91160 112534 91216
rect 112590 91160 112595 91216
rect 112364 91158 112595 91160
rect 112364 91156 112370 91158
rect 112529 91155 112595 91158
rect 113214 91156 113220 91220
rect 113284 91218 113290 91220
rect 114461 91218 114527 91221
rect 115841 91220 115907 91221
rect 117129 91220 117195 91221
rect 115790 91218 115796 91220
rect 113284 91216 114527 91218
rect 113284 91160 114466 91216
rect 114522 91160 114527 91216
rect 113284 91158 114527 91160
rect 115750 91158 115796 91218
rect 115860 91216 115907 91220
rect 117078 91218 117084 91220
rect 115902 91160 115907 91216
rect 113284 91156 113290 91158
rect 114461 91155 114527 91158
rect 115790 91156 115796 91158
rect 115860 91156 115907 91160
rect 117038 91158 117084 91218
rect 117148 91216 117195 91220
rect 117190 91160 117195 91216
rect 117078 91156 117084 91158
rect 117148 91156 117195 91160
rect 117998 91156 118004 91220
rect 118068 91218 118074 91220
rect 118601 91218 118667 91221
rect 118068 91216 118667 91218
rect 118068 91160 118606 91216
rect 118662 91160 118667 91216
rect 118068 91158 118667 91160
rect 118068 91156 118074 91158
rect 115841 91155 115907 91156
rect 117129 91155 117195 91156
rect 118601 91155 118667 91158
rect 119654 91156 119660 91220
rect 119724 91218 119730 91220
rect 119981 91218 120047 91221
rect 119724 91216 120047 91218
rect 119724 91160 119986 91216
rect 120042 91160 120047 91216
rect 119724 91158 120047 91160
rect 119724 91156 119730 91158
rect 119981 91155 120047 91158
rect 120206 91156 120212 91220
rect 120276 91218 120282 91220
rect 121361 91218 121427 91221
rect 120276 91216 121427 91218
rect 120276 91160 121366 91216
rect 121422 91160 121427 91216
rect 120276 91158 121427 91160
rect 120276 91156 120282 91158
rect 121361 91155 121427 91158
rect 122046 91156 122052 91220
rect 122116 91218 122122 91220
rect 122741 91218 122807 91221
rect 122116 91216 122807 91218
rect 122116 91160 122746 91216
rect 122802 91160 122807 91216
rect 122116 91158 122807 91160
rect 122116 91156 122122 91158
rect 122741 91155 122807 91158
rect 123150 91156 123156 91220
rect 123220 91218 123226 91220
rect 124121 91218 124187 91221
rect 123220 91216 124187 91218
rect 123220 91160 124126 91216
rect 124182 91160 124187 91216
rect 123220 91158 124187 91160
rect 123220 91156 123226 91158
rect 124121 91155 124187 91158
rect 125358 91156 125364 91220
rect 125428 91218 125434 91220
rect 125501 91218 125567 91221
rect 125428 91216 125567 91218
rect 125428 91160 125506 91216
rect 125562 91160 125567 91216
rect 125428 91158 125567 91160
rect 125428 91156 125434 91158
rect 125501 91155 125567 91158
rect 130694 91156 130700 91220
rect 130764 91218 130770 91220
rect 131021 91218 131087 91221
rect 132401 91220 132467 91221
rect 132350 91218 132356 91220
rect 130764 91216 131087 91218
rect 130764 91160 131026 91216
rect 131082 91160 131087 91216
rect 130764 91158 131087 91160
rect 132310 91158 132356 91218
rect 132420 91216 132467 91220
rect 132462 91160 132467 91216
rect 130764 91156 130770 91158
rect 131021 91155 131087 91158
rect 132350 91156 132356 91158
rect 132420 91156 132467 91160
rect 133086 91156 133092 91220
rect 133156 91218 133162 91220
rect 133229 91218 133295 91221
rect 133156 91216 133295 91218
rect 133156 91160 133234 91216
rect 133290 91160 133295 91216
rect 133156 91158 133295 91160
rect 133156 91156 133162 91158
rect 132401 91155 132467 91156
rect 133229 91155 133295 91158
rect 151486 91156 151492 91220
rect 151556 91218 151562 91220
rect 151721 91218 151787 91221
rect 151556 91216 151787 91218
rect 151556 91160 151726 91216
rect 151782 91160 151787 91216
rect 151556 91158 151787 91160
rect 151556 91156 151562 91158
rect 151721 91155 151787 91158
rect 168230 91082 168236 91084
rect 98134 91022 168236 91082
rect 168230 91020 168236 91022
rect 168300 91020 168306 91084
rect 106089 89722 106155 89725
rect 162853 89722 162919 89725
rect 106089 89720 162919 89722
rect 106089 89664 106094 89720
rect 106150 89664 162858 89720
rect 162914 89664 162919 89720
rect 106089 89662 162919 89664
rect 106089 89659 106155 89662
rect 162853 89659 162919 89662
rect 110689 88226 110755 88229
rect 166390 88226 166396 88228
rect 110689 88224 166396 88226
rect 110689 88168 110694 88224
rect 110750 88168 166396 88224
rect 110689 88166 166396 88168
rect 110689 88163 110755 88166
rect 166390 88164 166396 88166
rect 166460 88164 166466 88228
rect 88057 86866 88123 86869
rect 170254 86866 170260 86868
rect 88057 86864 170260 86866
rect 88057 86808 88062 86864
rect 88118 86808 170260 86864
rect 88057 86806 170260 86808
rect 88057 86803 88123 86806
rect 170254 86804 170260 86806
rect 170324 86804 170330 86868
rect 583017 86186 583083 86189
rect 583520 86186 584960 86276
rect 583017 86184 584960 86186
rect 583017 86128 583022 86184
rect 583078 86128 584960 86184
rect 583017 86126 584960 86128
rect 583017 86123 583083 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 103421 84146 103487 84149
rect 166206 84146 166212 84148
rect 103421 84144 166212 84146
rect 103421 84088 103426 84144
rect 103482 84088 166212 84144
rect 103421 84086 166212 84088
rect 103421 84083 103487 84086
rect 166206 84084 166212 84086
rect 166276 84084 166282 84148
rect 119889 84010 119955 84013
rect 170438 84010 170444 84012
rect 119889 84008 170444 84010
rect 119889 83952 119894 84008
rect 119950 83952 170444 84008
rect 119889 83950 170444 83952
rect 119889 83947 119955 83950
rect 170438 83948 170444 83950
rect 170508 83948 170514 84012
rect 66069 81426 66135 81429
rect 214414 81426 214420 81428
rect 66069 81424 214420 81426
rect 66069 81368 66074 81424
rect 66130 81368 214420 81424
rect 66069 81366 214420 81368
rect 66069 81363 66135 81366
rect 214414 81364 214420 81366
rect 214484 81364 214490 81428
rect 178534 80684 178540 80748
rect 178604 80746 178610 80748
rect 255313 80746 255379 80749
rect 178604 80744 255379 80746
rect 178604 80688 255318 80744
rect 255374 80688 255379 80744
rect 178604 80686 255379 80688
rect 178604 80684 178610 80686
rect 255313 80683 255379 80686
rect 99281 80066 99347 80069
rect 168966 80066 168972 80068
rect 99281 80064 168972 80066
rect 99281 80008 99286 80064
rect 99342 80008 168972 80064
rect 99281 80006 168972 80008
rect 99281 80003 99347 80006
rect 168966 80004 168972 80006
rect 169036 80004 169042 80068
rect 582465 72994 582531 72997
rect 583520 72994 584960 73084
rect 582465 72992 584960 72994
rect 582465 72936 582470 72992
rect 582526 72936 584960 72992
rect 582465 72934 584960 72936
rect 582465 72931 582531 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 56593 64154 56659 64157
rect 304206 64154 304212 64156
rect 56593 64152 304212 64154
rect 56593 64096 56598 64152
rect 56654 64096 304212 64152
rect 56593 64094 304212 64096
rect 56593 64091 56659 64094
rect 304206 64092 304212 64094
rect 304276 64092 304282 64156
rect 49693 62794 49759 62797
rect 305494 62794 305500 62796
rect 49693 62792 305500 62794
rect 49693 62736 49698 62792
rect 49754 62736 305500 62792
rect 49693 62734 305500 62736
rect 49693 62731 49759 62734
rect 305494 62732 305500 62734
rect 305564 62732 305570 62796
rect 582741 59666 582807 59669
rect 583520 59666 584960 59756
rect 582741 59664 584960 59666
rect 582741 59608 582746 59664
rect 582802 59608 584960 59664
rect 582741 59606 584960 59608
rect 582741 59603 582807 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 22093 53138 22159 53141
rect 299974 53138 299980 53140
rect 22093 53136 299980 53138
rect 22093 53080 22098 53136
rect 22154 53080 299980 53136
rect 22093 53078 299980 53080
rect 22093 53075 22159 53078
rect 299974 53076 299980 53078
rect 300044 53076 300050 53140
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 2773 36546 2839 36549
rect 302734 36546 302740 36548
rect 2773 36544 302740 36546
rect 2773 36488 2778 36544
rect 2834 36488 302740 36544
rect 2773 36486 302740 36488
rect 2773 36483 2839 36486
rect 302734 36484 302740 36486
rect 302804 36484 302810 36548
rect 271086 33764 271092 33828
rect 271156 33826 271162 33828
rect 296713 33826 296779 33829
rect 271156 33824 296779 33826
rect 271156 33768 296718 33824
rect 296774 33768 296779 33824
rect 271156 33766 296779 33768
rect 271156 33764 271162 33766
rect 296713 33763 296779 33766
rect 582833 33146 582899 33149
rect 583520 33146 584960 33236
rect 582833 33144 584960 33146
rect 582833 33088 582838 33144
rect 582894 33088 584960 33144
rect 582833 33086 584960 33088
rect 582833 33083 582899 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 64638 30908 64644 30972
rect 64708 30970 64714 30972
rect 307845 30970 307911 30973
rect 64708 30968 307911 30970
rect 64708 30912 307850 30968
rect 307906 30912 307911 30968
rect 64708 30910 307911 30912
rect 64708 30908 64714 30910
rect 307845 30907 307911 30910
rect 62982 26828 62988 26892
rect 63052 26890 63058 26892
rect 248413 26890 248479 26893
rect 63052 26888 248479 26890
rect 63052 26832 248418 26888
rect 248474 26832 248479 26888
rect 63052 26830 248479 26832
rect 63052 26828 63058 26830
rect 248413 26827 248479 26830
rect 77385 19954 77451 19957
rect 253054 19954 253060 19956
rect 77385 19952 253060 19954
rect 77385 19896 77390 19952
rect 77446 19896 253060 19952
rect 77385 19894 253060 19896
rect 77385 19891 77451 19894
rect 253054 19892 253060 19894
rect 253124 19892 253130 19956
rect 582373 19818 582439 19821
rect 583520 19818 584960 19908
rect 582373 19816 584960 19818
rect 582373 19760 582378 19816
rect 582434 19760 584960 19816
rect 582373 19758 584960 19760
rect 582373 19755 582439 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 269614 14452 269620 14516
rect 269684 14514 269690 14516
rect 299473 14514 299539 14517
rect 269684 14512 299539 14514
rect 269684 14456 299478 14512
rect 299534 14456 299539 14512
rect 269684 14454 299539 14456
rect 269684 14452 269690 14454
rect 299473 14451 299539 14454
rect 66110 13092 66116 13156
rect 66180 13154 66186 13156
rect 251265 13154 251331 13157
rect 66180 13152 251331 13154
rect 66180 13096 251270 13152
rect 251326 13096 251331 13152
rect 66180 13094 251331 13096
rect 66180 13092 66186 13094
rect 251265 13091 251331 13094
rect 9673 13018 9739 13021
rect 306966 13018 306972 13020
rect 9673 13016 306972 13018
rect 9673 12960 9678 13016
rect 9734 12960 306972 13016
rect 9673 12958 306972 12960
rect 9673 12955 9739 12958
rect 306966 12956 306972 12958
rect 307036 12956 307042 13020
rect 582649 6626 582715 6629
rect 583520 6626 584960 6716
rect 582649 6624 584960 6626
rect -960 6490 480 6580
rect 582649 6568 582654 6624
rect 582710 6568 584960 6624
rect 582649 6566 584960 6568
rect 582649 6563 582715 6566
rect 4061 6490 4127 6493
rect -960 6488 4127 6490
rect -960 6432 4066 6488
rect 4122 6432 4127 6488
rect 583520 6476 584960 6566
rect -960 6430 4127 6432
rect -960 6340 480 6430
rect 4061 6427 4127 6430
rect 15193 4858 15259 4861
rect 307150 4858 307156 4860
rect 15193 4856 307156 4858
rect 15193 4800 15198 4856
rect 15254 4800 307156 4856
rect 15193 4798 307156 4800
rect 15193 4795 15259 4798
rect 307150 4796 307156 4798
rect 307220 4796 307226 4860
rect 335118 3980 335124 4044
rect 335188 4042 335194 4044
rect 336273 4042 336339 4045
rect 335188 4040 336339 4042
rect 335188 3984 336278 4040
rect 336334 3984 336339 4040
rect 335188 3982 336339 3984
rect 335188 3980 335194 3982
rect 336273 3979 336339 3982
rect 262806 3572 262812 3636
rect 262876 3634 262882 3636
rect 262876 3574 266738 3634
rect 262876 3572 262882 3574
rect 258257 3498 258323 3501
rect 259453 3500 259519 3501
rect 258390 3498 258396 3500
rect 258257 3496 258396 3498
rect 258257 3440 258262 3496
rect 258318 3440 258396 3496
rect 258257 3438 258396 3440
rect 258257 3435 258323 3438
rect 258390 3436 258396 3438
rect 258460 3436 258466 3500
rect 259453 3498 259500 3500
rect 259408 3496 259500 3498
rect 259408 3440 259458 3496
rect 259408 3438 259500 3440
rect 259453 3436 259500 3438
rect 259564 3436 259570 3500
rect 263542 3436 263548 3500
rect 263612 3498 263618 3500
rect 264145 3498 264211 3501
rect 263612 3496 264211 3498
rect 263612 3440 264150 3496
rect 264206 3440 264211 3496
rect 263612 3438 264211 3440
rect 263612 3436 263618 3438
rect 259453 3435 259519 3436
rect 264145 3435 264211 3438
rect 265341 3498 265407 3501
rect 265750 3498 265756 3500
rect 265341 3496 265756 3498
rect 265341 3440 265346 3496
rect 265402 3440 265756 3496
rect 265341 3438 265756 3440
rect 265341 3435 265407 3438
rect 265750 3436 265756 3438
rect 265820 3436 265826 3500
rect 266302 3436 266308 3500
rect 266372 3498 266378 3500
rect 266537 3498 266603 3501
rect 266372 3496 266603 3498
rect 266372 3440 266542 3496
rect 266598 3440 266603 3496
rect 266372 3438 266603 3440
rect 266678 3498 266738 3574
rect 267774 3572 267780 3636
rect 267844 3634 267850 3636
rect 268837 3634 268903 3637
rect 267844 3632 268903 3634
rect 267844 3576 268842 3632
rect 268898 3576 268903 3632
rect 267844 3574 268903 3576
rect 267844 3572 267850 3574
rect 268837 3571 268903 3574
rect 276238 3572 276244 3636
rect 276308 3634 276314 3636
rect 277117 3634 277183 3637
rect 276308 3632 277183 3634
rect 276308 3576 277122 3632
rect 277178 3576 277183 3632
rect 276308 3574 277183 3576
rect 276308 3572 276314 3574
rect 277117 3571 277183 3574
rect 286174 3572 286180 3636
rect 286244 3634 286250 3636
rect 290181 3634 290247 3637
rect 286244 3632 290247 3634
rect 286244 3576 290186 3632
rect 290242 3576 290247 3632
rect 286244 3574 290247 3576
rect 286244 3572 286250 3574
rect 290181 3571 290247 3574
rect 298686 3572 298692 3636
rect 298756 3634 298762 3636
rect 298756 3574 306390 3634
rect 298756 3572 298762 3574
rect 286593 3498 286659 3501
rect 266678 3496 286659 3498
rect 266678 3440 286598 3496
rect 286654 3440 286659 3496
rect 266678 3438 286659 3440
rect 266372 3436 266378 3438
rect 266537 3435 266603 3438
rect 286593 3435 286659 3438
rect 288382 3436 288388 3500
rect 288452 3498 288458 3500
rect 288985 3498 289051 3501
rect 288452 3496 289051 3498
rect 288452 3440 288990 3496
rect 289046 3440 289051 3496
rect 288452 3438 289051 3440
rect 288452 3436 288458 3438
rect 288985 3435 289051 3438
rect 301814 3436 301820 3500
rect 301884 3498 301890 3500
rect 301957 3498 302023 3501
rect 301884 3496 302023 3498
rect 301884 3440 301962 3496
rect 302018 3440 302023 3496
rect 301884 3438 302023 3440
rect 301884 3436 301890 3438
rect 301957 3435 302023 3438
rect 302182 3436 302188 3500
rect 302252 3498 302258 3500
rect 303153 3498 303219 3501
rect 302252 3496 303219 3498
rect 302252 3440 303158 3496
rect 303214 3440 303219 3496
rect 302252 3438 303219 3440
rect 302252 3436 302258 3438
rect 303153 3435 303219 3438
rect 303654 3436 303660 3500
rect 303724 3498 303730 3500
rect 304349 3498 304415 3501
rect 303724 3496 304415 3498
rect 303724 3440 304354 3496
rect 304410 3440 304415 3496
rect 303724 3438 304415 3440
rect 303724 3436 303730 3438
rect 304349 3435 304415 3438
rect 304942 3436 304948 3500
rect 305012 3498 305018 3500
rect 305545 3498 305611 3501
rect 305012 3496 305611 3498
rect 305012 3440 305550 3496
rect 305606 3440 305611 3496
rect 305012 3438 305611 3440
rect 306330 3498 306390 3574
rect 334014 3572 334020 3636
rect 334084 3634 334090 3636
rect 335077 3634 335143 3637
rect 334084 3632 335143 3634
rect 334084 3576 335082 3632
rect 335138 3576 335143 3632
rect 334084 3574 335143 3576
rect 334084 3572 334090 3574
rect 335077 3571 335143 3574
rect 319713 3498 319779 3501
rect 306330 3496 319779 3498
rect 306330 3440 319718 3496
rect 319774 3440 319779 3496
rect 306330 3438 319779 3440
rect 305012 3436 305018 3438
rect 305545 3435 305611 3438
rect 319713 3435 319779 3438
rect 331254 3436 331260 3500
rect 331324 3498 331330 3500
rect 331581 3498 331647 3501
rect 331324 3496 331647 3498
rect 331324 3440 331586 3496
rect 331642 3440 331647 3496
rect 331324 3438 331647 3440
rect 331324 3436 331330 3438
rect 331581 3435 331647 3438
rect 332542 3436 332548 3500
rect 332612 3498 332618 3500
rect 332685 3498 332751 3501
rect 332612 3496 332751 3498
rect 332612 3440 332690 3496
rect 332746 3440 332751 3496
rect 332612 3438 332751 3440
rect 332612 3436 332618 3438
rect 332685 3435 332751 3438
rect 333881 3498 333947 3501
rect 334198 3498 334204 3500
rect 333881 3496 334204 3498
rect 333881 3440 333886 3496
rect 333942 3440 334204 3496
rect 333881 3438 334204 3440
rect 333881 3435 333947 3438
rect 334198 3436 334204 3438
rect 334268 3436 334274 3500
rect 335854 3436 335860 3500
rect 335924 3498 335930 3500
rect 337469 3498 337535 3501
rect 335924 3496 337535 3498
rect 335924 3440 337474 3496
rect 337530 3440 337535 3496
rect 335924 3438 337535 3440
rect 335924 3436 335930 3438
rect 337469 3435 337535 3438
rect 338246 3436 338252 3500
rect 338316 3498 338322 3500
rect 338665 3498 338731 3501
rect 338316 3496 338731 3498
rect 338316 3440 338670 3496
rect 338726 3440 338731 3496
rect 338316 3438 338731 3440
rect 338316 3436 338322 3438
rect 338665 3435 338731 3438
rect 339534 3436 339540 3500
rect 339604 3498 339610 3500
rect 339861 3498 339927 3501
rect 339604 3496 339927 3498
rect 339604 3440 339866 3496
rect 339922 3440 339927 3496
rect 339604 3438 339927 3440
rect 339604 3436 339610 3438
rect 339861 3435 339927 3438
rect 340822 3436 340828 3500
rect 340892 3498 340898 3500
rect 340965 3498 341031 3501
rect 340892 3496 341031 3498
rect 340892 3440 340970 3496
rect 341026 3440 341031 3496
rect 340892 3438 341031 3440
rect 340892 3436 340898 3438
rect 340965 3435 341031 3438
rect 342294 3436 342300 3500
rect 342364 3498 342370 3500
rect 343357 3498 343423 3501
rect 342364 3496 343423 3498
rect 342364 3440 343362 3496
rect 343418 3440 343423 3496
rect 342364 3438 343423 3440
rect 342364 3436 342370 3438
rect 343357 3435 343423 3438
rect 345054 3436 345060 3500
rect 345124 3498 345130 3500
rect 345749 3498 345815 3501
rect 345124 3496 345815 3498
rect 345124 3440 345754 3496
rect 345810 3440 345815 3496
rect 345124 3438 345815 3440
rect 345124 3436 345130 3438
rect 345749 3435 345815 3438
rect 273846 3300 273852 3364
rect 273916 3362 273922 3364
rect 299657 3362 299723 3365
rect 273916 3360 299723 3362
rect 273916 3304 299662 3360
rect 299718 3304 299723 3360
rect 273916 3302 299723 3304
rect 273916 3300 273922 3302
rect 299657 3299 299723 3302
<< via3 >>
rect 69060 696900 69124 696964
rect 177252 387772 177316 387836
rect 57836 383828 57900 383892
rect 273852 383692 273916 383756
rect 170260 381244 170324 381308
rect 262812 381108 262876 381172
rect 286180 380972 286244 381036
rect 303660 380156 303724 380220
rect 298692 379476 298756 379540
rect 259500 379068 259564 379132
rect 304948 377708 305012 377772
rect 109356 377028 109420 377092
rect 178540 373628 178604 373692
rect 110644 373356 110708 373420
rect 65932 370228 65996 370292
rect 269620 368460 269684 368524
rect 66668 366148 66732 366212
rect 335860 366284 335924 366348
rect 267780 364924 267844 364988
rect 64644 360300 64708 360364
rect 276244 357988 276308 358052
rect 271092 353500 271156 353564
rect 301820 352548 301884 352612
rect 66116 347108 66180 347172
rect 62988 346564 63052 346628
rect 125732 343708 125796 343772
rect 69060 343572 69124 343636
rect 70348 343028 70412 343092
rect 331260 340036 331324 340100
rect 65932 339900 65996 339964
rect 124260 339356 124324 339420
rect 61884 337452 61948 337516
rect 70348 337316 70412 337380
rect 108988 336636 109052 336700
rect 58940 335956 59004 336020
rect 266308 334596 266372 334660
rect 59124 333236 59188 333300
rect 118740 331876 118804 331940
rect 66668 331740 66732 331804
rect 338252 331740 338316 331804
rect 263548 330380 263612 330444
rect 339540 327660 339604 327724
rect 288388 325076 288452 325140
rect 342300 324940 342364 325004
rect 340828 319364 340892 319428
rect 265756 313924 265820 313988
rect 345060 309708 345124 309772
rect 302188 305628 302252 305692
rect 334020 304132 334084 304196
rect 70900 301548 70964 301612
rect 258396 301412 258460 301476
rect 110644 300052 110708 300116
rect 321508 296788 321572 296852
rect 252508 295428 252572 295492
rect 123340 294204 123404 294268
rect 322980 293932 323044 293996
rect 327028 291892 327092 291956
rect 65932 289172 65996 289236
rect 70532 286724 70596 286788
rect 123340 282100 123404 282164
rect 580212 282100 580276 282164
rect 255268 274620 255332 274684
rect 61700 254008 61764 254012
rect 61700 253952 61714 254008
rect 61714 253952 61764 254008
rect 61700 253948 61764 253952
rect 332548 253132 332612 253196
rect 58940 245652 59004 245716
rect 59124 241708 59188 241772
rect 57836 240348 57900 240412
rect 119292 240892 119356 240956
rect 118740 239804 118804 239868
rect 125732 238580 125796 238644
rect 124260 238444 124324 238508
rect 61884 237220 61948 237284
rect 61700 232460 61764 232524
rect 328500 226884 328564 226948
rect 258396 218588 258460 218652
rect 65932 217228 65996 217292
rect 262260 211788 262324 211852
rect 336780 206212 336844 206276
rect 118924 200636 118988 200700
rect 339724 192476 339788 192540
rect 259684 186900 259748 186964
rect 256740 185540 256804 185604
rect 331444 180100 331508 180164
rect 338252 179964 338316 180028
rect 166212 179420 166276 179484
rect 266492 178740 266556 178804
rect 98316 177652 98380 177716
rect 104572 177652 104636 177716
rect 106964 177652 107028 177716
rect 110644 177712 110708 177716
rect 110644 177656 110694 177712
rect 110694 177656 110708 177712
rect 110644 177652 110708 177656
rect 114324 177652 114388 177716
rect 115796 177712 115860 177716
rect 115796 177656 115846 177712
rect 115846 177656 115860 177712
rect 115796 177652 115860 177656
rect 116900 177712 116964 177716
rect 116900 177656 116950 177712
rect 116950 177656 116964 177712
rect 116900 177652 116964 177656
rect 119476 177652 119540 177716
rect 120764 177652 120828 177716
rect 129412 177652 129476 177716
rect 130700 177712 130764 177716
rect 130700 177656 130750 177712
rect 130750 177656 130764 177712
rect 130700 177652 130764 177656
rect 249196 177516 249260 177580
rect 249380 177380 249444 177444
rect 335124 177380 335188 177444
rect 334204 177244 334268 177308
rect 97028 176972 97092 177036
rect 112116 177032 112180 177036
rect 112116 176976 112166 177032
rect 112166 176976 112180 177032
rect 112116 176972 112180 176976
rect 124444 176972 124508 177036
rect 105676 176836 105740 176900
rect 168236 176836 168300 176900
rect 101996 176760 102060 176764
rect 101996 176704 102046 176760
rect 102046 176704 102060 176760
rect 101996 176700 102060 176704
rect 108068 176760 108132 176764
rect 108068 176704 108118 176760
rect 108118 176704 108132 176760
rect 108068 176700 108132 176704
rect 109540 176700 109604 176764
rect 123156 176700 123220 176764
rect 125732 176700 125796 176764
rect 133092 176760 133156 176764
rect 133092 176704 133142 176760
rect 133142 176704 133156 176760
rect 133092 176700 133156 176704
rect 134380 176760 134444 176764
rect 134380 176704 134430 176760
rect 134430 176704 134444 176760
rect 134380 176700 134444 176704
rect 136036 176760 136100 176764
rect 136036 176704 136086 176760
rect 136086 176704 136100 176760
rect 136036 176700 136100 176704
rect 148180 176760 148244 176764
rect 148180 176704 148230 176760
rect 148230 176704 148244 176760
rect 148180 176700 148244 176704
rect 99420 176428 99484 176492
rect 103284 176428 103348 176492
rect 128124 176428 128188 176492
rect 263732 176292 263796 176356
rect 113220 175476 113284 175540
rect 127020 175536 127084 175540
rect 127020 175480 127070 175536
rect 127070 175480 127084 175536
rect 100708 175400 100772 175404
rect 100708 175344 100758 175400
rect 100758 175344 100772 175400
rect 100708 175340 100772 175344
rect 118372 175400 118436 175404
rect 118372 175344 118422 175400
rect 118422 175344 118436 175400
rect 118372 175340 118436 175344
rect 121868 175400 121932 175404
rect 121868 175344 121918 175400
rect 121918 175344 121932 175400
rect 121868 175340 121932 175344
rect 127020 175476 127084 175480
rect 131988 175536 132052 175540
rect 131988 175480 132038 175536
rect 132038 175480 132052 175536
rect 131988 175476 132052 175480
rect 158852 175536 158916 175540
rect 158852 175480 158902 175536
rect 158902 175480 158916 175536
rect 158852 175476 158916 175480
rect 166396 175340 166460 175404
rect 262076 175340 262140 175404
rect 306972 175204 307036 175268
rect 249196 174660 249260 174724
rect 249380 173300 249444 173364
rect 166396 163100 166460 163164
rect 262260 161740 262324 161804
rect 258396 159292 258460 159356
rect 168236 158748 168300 158812
rect 259684 158612 259748 158676
rect 263732 157116 263796 157180
rect 166212 154532 166276 154596
rect 255268 152084 255332 152148
rect 256740 147460 256804 147524
rect 251772 142700 251836 142764
rect 254532 141476 254596 141540
rect 306972 141340 307036 141404
rect 307524 141204 307588 141268
rect 266492 141068 266556 141132
rect 302740 139708 302804 139772
rect 580212 139300 580276 139364
rect 170444 138076 170508 138140
rect 252508 137940 252572 138004
rect 169156 135220 169220 135284
rect 166396 134132 166460 134196
rect 321508 134404 321572 134468
rect 253060 134132 253124 134196
rect 307524 131684 307588 131748
rect 327028 131684 327092 131748
rect 304212 131412 304276 131476
rect 166212 130052 166276 130116
rect 305500 130052 305564 130116
rect 168972 128556 169036 128620
rect 168236 127060 168300 127124
rect 306972 126380 307036 126444
rect 339724 124204 339788 124268
rect 336780 115908 336844 115972
rect 170260 115092 170324 115156
rect 299980 113868 300044 113932
rect 331444 111012 331508 111076
rect 322980 107068 323044 107132
rect 177252 106796 177316 106860
rect 328500 106252 328564 106316
rect 173020 105164 173084 105228
rect 214604 105028 214668 105092
rect 251772 104620 251836 104684
rect 254532 101764 254596 101828
rect 338252 100948 338316 101012
rect 170260 99452 170324 99516
rect 214420 97004 214484 97068
rect 307156 97004 307220 97068
rect 324452 97004 324516 97068
rect 262076 96596 262140 96660
rect 173020 94828 173084 94892
rect 106228 94692 106292 94756
rect 106614 94692 106678 94756
rect 129326 94752 129390 94756
rect 129326 94696 129370 94752
rect 129370 94696 129390 94752
rect 129326 94692 129390 94696
rect 151766 94752 151830 94756
rect 151766 94696 151782 94752
rect 151782 94696 151830 94752
rect 151766 94692 151830 94696
rect 111932 93876 111996 93940
rect 169156 93876 169220 93940
rect 214604 93740 214668 93804
rect 85620 93664 85684 93668
rect 85620 93608 85670 93664
rect 85670 93608 85684 93664
rect 85620 93604 85684 93608
rect 115428 93664 115492 93668
rect 115428 93608 115478 93664
rect 115478 93608 115492 93664
rect 115428 93604 115492 93608
rect 120580 93664 120644 93668
rect 120580 93608 120630 93664
rect 120630 93608 120644 93664
rect 120580 93604 120644 93608
rect 135668 93664 135732 93668
rect 135668 93608 135718 93664
rect 135718 93608 135732 93664
rect 135668 93604 135732 93608
rect 151676 93664 151740 93668
rect 151676 93608 151726 93664
rect 151726 93608 151740 93664
rect 151676 93604 151740 93608
rect 324452 93604 324516 93668
rect 103284 93196 103348 93260
rect 110276 93256 110340 93260
rect 110276 93200 110326 93256
rect 110326 93200 110340 93256
rect 110276 93196 110340 93200
rect 113772 93256 113836 93260
rect 113772 93200 113822 93256
rect 113822 93200 113836 93256
rect 113772 93196 113836 93200
rect 128124 93256 128188 93260
rect 128124 93200 128174 93256
rect 128174 93200 128188 93256
rect 128124 93196 128188 93200
rect 74764 92440 74828 92444
rect 74764 92384 74814 92440
rect 74814 92384 74828 92440
rect 74764 92380 74828 92384
rect 88932 92440 88996 92444
rect 88932 92384 88982 92440
rect 88982 92384 88996 92440
rect 88932 92380 88996 92384
rect 95004 92440 95068 92444
rect 95004 92384 95054 92440
rect 95054 92384 95068 92440
rect 95004 92380 95068 92384
rect 101812 92380 101876 92444
rect 105492 92440 105556 92444
rect 105492 92384 105542 92440
rect 105542 92384 105556 92440
rect 105492 92380 105556 92384
rect 106228 92380 106292 92444
rect 116716 92440 116780 92444
rect 116716 92384 116766 92440
rect 116766 92384 116780 92440
rect 116716 92380 116780 92384
rect 124076 92440 124140 92444
rect 124076 92384 124090 92440
rect 124090 92384 124140 92440
rect 124076 92380 124140 92384
rect 125732 92380 125796 92444
rect 134380 92440 134444 92444
rect 134380 92384 134430 92440
rect 134430 92384 134444 92440
rect 134380 92380 134444 92384
rect 152044 92380 152108 92444
rect 114324 92244 114388 92308
rect 126652 92032 126716 92036
rect 126652 91976 126702 92032
rect 126702 91976 126716 92032
rect 126652 91972 126716 91976
rect 105676 91700 105740 91764
rect 114876 91700 114940 91764
rect 124444 91564 124508 91628
rect 126468 91564 126532 91628
rect 122788 91488 122852 91492
rect 122788 91432 122838 91488
rect 122838 91432 122852 91488
rect 122788 91428 122852 91432
rect 98500 91292 98564 91356
rect 100892 91292 100956 91356
rect 104204 91292 104268 91356
rect 108068 91292 108132 91356
rect 109540 91352 109604 91356
rect 109540 91296 109590 91352
rect 109590 91296 109604 91352
rect 109540 91292 109604 91296
rect 118188 91352 118252 91356
rect 118188 91296 118238 91352
rect 118238 91296 118252 91352
rect 118188 91292 118252 91296
rect 119292 91292 119356 91356
rect 121684 91292 121748 91356
rect 84332 91156 84396 91220
rect 86724 91156 86788 91220
rect 88012 91216 88076 91220
rect 88012 91160 88062 91216
rect 88062 91160 88076 91216
rect 88012 91156 88076 91160
rect 90220 91156 90284 91220
rect 91324 91156 91388 91220
rect 92612 91156 92676 91220
rect 93900 91156 93964 91220
rect 96292 91156 96356 91220
rect 96660 91156 96724 91220
rect 97212 91156 97276 91220
rect 98132 91156 98196 91220
rect 99052 91156 99116 91220
rect 99972 91156 100036 91220
rect 100524 91156 100588 91220
rect 101996 91216 102060 91220
rect 101996 91160 102010 91216
rect 102010 91160 102060 91216
rect 101996 91156 102060 91160
rect 102732 91156 102796 91220
rect 104572 91156 104636 91220
rect 106596 91156 106660 91220
rect 107700 91156 107764 91220
rect 109172 91156 109236 91220
rect 110644 91216 110708 91220
rect 110644 91160 110694 91216
rect 110694 91160 110708 91216
rect 110644 91156 110708 91160
rect 111196 91156 111260 91220
rect 112300 91156 112364 91220
rect 113220 91156 113284 91220
rect 115796 91216 115860 91220
rect 115796 91160 115846 91216
rect 115846 91160 115860 91216
rect 115796 91156 115860 91160
rect 117084 91216 117148 91220
rect 117084 91160 117134 91216
rect 117134 91160 117148 91216
rect 117084 91156 117148 91160
rect 118004 91156 118068 91220
rect 119660 91156 119724 91220
rect 120212 91156 120276 91220
rect 122052 91156 122116 91220
rect 123156 91156 123220 91220
rect 125364 91156 125428 91220
rect 130700 91156 130764 91220
rect 132356 91216 132420 91220
rect 132356 91160 132406 91216
rect 132406 91160 132420 91216
rect 132356 91156 132420 91160
rect 133092 91156 133156 91220
rect 151492 91156 151556 91220
rect 168236 91020 168300 91084
rect 166396 88164 166460 88228
rect 170260 86804 170324 86868
rect 166212 84084 166276 84148
rect 170444 83948 170508 84012
rect 214420 81364 214484 81428
rect 178540 80684 178604 80748
rect 168972 80004 169036 80068
rect 304212 64092 304276 64156
rect 305500 62732 305564 62796
rect 299980 53076 300044 53140
rect 302740 36484 302804 36548
rect 271092 33764 271156 33828
rect 64644 30908 64708 30972
rect 62988 26828 63052 26892
rect 253060 19892 253124 19956
rect 269620 14452 269684 14516
rect 66116 13092 66180 13156
rect 306972 12956 307036 13020
rect 307156 4796 307220 4860
rect 335124 3980 335188 4044
rect 262812 3572 262876 3636
rect 258396 3436 258460 3500
rect 259500 3496 259564 3500
rect 259500 3440 259514 3496
rect 259514 3440 259564 3496
rect 259500 3436 259564 3440
rect 263548 3436 263612 3500
rect 265756 3436 265820 3500
rect 266308 3436 266372 3500
rect 267780 3572 267844 3636
rect 276244 3572 276308 3636
rect 286180 3572 286244 3636
rect 298692 3572 298756 3636
rect 288388 3436 288452 3500
rect 301820 3436 301884 3500
rect 302188 3436 302252 3500
rect 303660 3436 303724 3500
rect 304948 3436 305012 3500
rect 334020 3572 334084 3636
rect 331260 3436 331324 3500
rect 332548 3436 332612 3500
rect 334204 3436 334268 3500
rect 335860 3436 335924 3500
rect 338252 3436 338316 3500
rect 339540 3436 339604 3500
rect 340828 3436 340892 3500
rect 342300 3436 342364 3500
rect 345060 3436 345124 3500
rect 273852 3300 273916 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 57835 383892 57901 383893
rect 57835 383828 57836 383892
rect 57900 383828 57901 383892
rect 57835 383827 57901 383828
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 57838 240413 57898 383827
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 58939 336020 59005 336021
rect 58939 335956 58940 336020
rect 59004 335956 59005 336020
rect 58939 335955 59005 335956
rect 58942 245717 59002 335955
rect 59123 333300 59189 333301
rect 59123 333236 59124 333300
rect 59188 333236 59189 333300
rect 59123 333235 59189 333236
rect 58939 245716 59005 245717
rect 58939 245652 58940 245716
rect 59004 245652 59005 245716
rect 58939 245651 59005 245652
rect 59126 241773 59186 333235
rect 59514 313174 60134 348618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 69059 696964 69125 696965
rect 69059 696900 69060 696964
rect 69124 696900 69125 696964
rect 69059 696899 69125 696900
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 65931 370292 65997 370293
rect 65931 370228 65932 370292
rect 65996 370228 65997 370292
rect 65931 370227 65997 370228
rect 64643 360364 64709 360365
rect 64643 360300 64644 360364
rect 64708 360300 64709 360364
rect 64643 360299 64709 360300
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 62987 346628 63053 346629
rect 62987 346564 62988 346628
rect 63052 346564 63053 346628
rect 62987 346563 63053 346564
rect 61883 337516 61949 337517
rect 61883 337452 61884 337516
rect 61948 337452 61949 337516
rect 61883 337451 61949 337452
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59123 241772 59189 241773
rect 59123 241708 59124 241772
rect 59188 241708 59189 241772
rect 59123 241707 59189 241708
rect 59514 241174 60134 276618
rect 61699 254012 61765 254013
rect 61699 253948 61700 254012
rect 61764 253948 61765 254012
rect 61699 253947 61765 253948
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 57835 240412 57901 240413
rect 57835 240348 57836 240412
rect 57900 240348 57901 240412
rect 57835 240347 57901 240348
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 205174 60134 240618
rect 61702 232525 61762 253947
rect 61886 237285 61946 337451
rect 61883 237284 61949 237285
rect 61883 237220 61884 237284
rect 61948 237220 61949 237284
rect 61883 237219 61949 237220
rect 61699 232524 61765 232525
rect 61699 232460 61700 232524
rect 61764 232460 61765 232524
rect 61699 232459 61765 232460
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 62990 26893 63050 346563
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 64646 30973 64706 360299
rect 65934 339965 65994 370227
rect 66667 366212 66733 366213
rect 66667 366148 66668 366212
rect 66732 366148 66733 366212
rect 66667 366147 66733 366148
rect 66115 347172 66181 347173
rect 66115 347108 66116 347172
rect 66180 347108 66181 347172
rect 66115 347107 66181 347108
rect 65931 339964 65997 339965
rect 65931 339900 65932 339964
rect 65996 339900 65997 339964
rect 65931 339899 65997 339900
rect 65931 289236 65997 289237
rect 65931 289172 65932 289236
rect 65996 289172 65997 289236
rect 65931 289171 65997 289172
rect 65934 217293 65994 289171
rect 65931 217292 65997 217293
rect 65931 217228 65932 217292
rect 65996 217228 65997 217292
rect 65931 217227 65997 217228
rect 64643 30972 64709 30973
rect 64643 30908 64644 30972
rect 64708 30908 64709 30972
rect 64643 30907 64709 30908
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 62987 26892 63053 26893
rect 62987 26828 62988 26892
rect 63052 26828 63053 26892
rect 62987 26827 63053 26828
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 -5146 63854 28338
rect 66118 13157 66178 347107
rect 66670 331805 66730 366147
rect 66954 356614 67574 392058
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66667 331804 66733 331805
rect 66667 331740 66668 331804
rect 66732 331740 66733 331804
rect 66667 331739 66733 331740
rect 66954 320614 67574 356058
rect 69062 343637 69122 696899
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 382000 74414 398898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 382000 78134 402618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 382000 81854 406338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 382000 85574 410058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 382000 92414 416898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 385174 96134 420618
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 382000 96134 384618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 424894 99854 460338
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 388894 99854 424338
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 382000 99854 388338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 382000 103574 392058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 382000 110414 398898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 109355 377092 109421 377093
rect 109355 377028 109356 377092
rect 109420 377028 109421 377092
rect 109355 377027 109421 377028
rect 109358 374010 109418 377027
rect 108990 373950 109418 374010
rect 74208 363454 74528 363486
rect 74208 363218 74250 363454
rect 74486 363218 74528 363454
rect 74208 363134 74528 363218
rect 74208 362898 74250 363134
rect 74486 362898 74528 363134
rect 74208 362866 74528 362898
rect 104928 363454 105248 363486
rect 104928 363218 104970 363454
rect 105206 363218 105248 363454
rect 104928 363134 105248 363218
rect 104928 362898 104970 363134
rect 105206 362898 105248 363134
rect 104928 362866 105248 362898
rect 89568 345454 89888 345486
rect 89568 345218 89610 345454
rect 89846 345218 89888 345454
rect 89568 345134 89888 345218
rect 89568 344898 89610 345134
rect 89846 344898 89888 345134
rect 89568 344866 89888 344898
rect 69059 343636 69125 343637
rect 69059 343572 69060 343636
rect 69124 343572 69125 343636
rect 69059 343571 69125 343572
rect 70347 343092 70413 343093
rect 70347 343028 70348 343092
rect 70412 343028 70413 343092
rect 70347 343027 70413 343028
rect 70350 337381 70410 343027
rect 70347 337380 70413 337381
rect 70347 337316 70348 337380
rect 70412 337316 70413 337380
rect 70347 337315 70413 337316
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 73794 327454 74414 338000
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 70899 301612 70965 301613
rect 70899 301548 70900 301612
rect 70964 301548 70965 301612
rect 70899 301547 70965 301548
rect 70902 287070 70962 301547
rect 73794 294000 74414 326898
rect 77514 331174 78134 338000
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 294000 78134 294618
rect 81234 334894 81854 338000
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 294000 81854 298338
rect 84954 302614 85574 338000
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 294000 85574 302058
rect 91794 309454 92414 338000
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 294000 92414 308898
rect 95514 313174 96134 338000
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 294000 96134 312618
rect 99234 316894 99854 338000
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 294000 99854 316338
rect 102954 320614 103574 338000
rect 108990 336701 109050 373950
rect 110643 373420 110709 373421
rect 110643 373356 110644 373420
rect 110708 373356 110709 373420
rect 110643 373355 110709 373356
rect 108987 336700 109053 336701
rect 108987 336636 108988 336700
rect 109052 336636 109053 336700
rect 108987 336635 109053 336636
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 294000 103574 320058
rect 109794 327454 110414 338000
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 294000 110414 326898
rect 110646 300117 110706 373355
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 110643 300116 110709 300117
rect 110643 300052 110644 300116
rect 110708 300052 110709 300116
rect 110643 300051 110709 300052
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 294000 114134 294618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 125731 343772 125797 343773
rect 125731 343708 125732 343772
rect 125796 343708 125797 343772
rect 125731 343707 125797 343708
rect 124259 339420 124325 339421
rect 124259 339356 124260 339420
rect 124324 339356 124325 339420
rect 124259 339355 124325 339356
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 118739 331940 118805 331941
rect 118739 331876 118740 331940
rect 118804 331876 118805 331940
rect 118739 331875 118805 331876
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 294000 117854 298338
rect 70534 287010 70962 287070
rect 70534 286789 70594 287010
rect 70531 286788 70597 286789
rect 70531 286724 70532 286788
rect 70596 286724 70597 286788
rect 70531 286723 70597 286724
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 89568 273454 89888 273486
rect 89568 273218 89610 273454
rect 89846 273218 89888 273454
rect 89568 273134 89888 273218
rect 89568 272898 89610 273134
rect 89846 272898 89888 273134
rect 89568 272866 89888 272898
rect 74208 255454 74528 255486
rect 74208 255218 74250 255454
rect 74486 255218 74528 255454
rect 74208 255134 74528 255218
rect 74208 254898 74250 255134
rect 74486 254898 74528 255134
rect 74208 254866 74528 254898
rect 104928 255454 105248 255486
rect 104928 255218 104970 255454
rect 105206 255218 105248 255454
rect 104928 255134 105248 255218
rect 104928 254898 104970 255134
rect 105206 254898 105248 255134
rect 104928 254866 105248 254898
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 118742 239869 118802 331875
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 294000 121574 302058
rect 123339 294268 123405 294269
rect 123339 294204 123340 294268
rect 123404 294204 123405 294268
rect 123339 294203 123405 294204
rect 123342 282165 123402 294203
rect 123339 282164 123405 282165
rect 123339 282100 123340 282164
rect 123404 282100 123405 282164
rect 123339 282099 123405 282100
rect 119291 240956 119357 240957
rect 119291 240892 119292 240956
rect 119356 240892 119357 240956
rect 119291 240891 119357 240892
rect 118739 239868 118805 239869
rect 118739 239804 118740 239868
rect 118804 239804 118805 239868
rect 118739 239803 118805 239804
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176600 67574 212058
rect 73794 219454 74414 238000
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 176600 74414 182898
rect 77514 223174 78134 238000
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 176600 78134 186618
rect 81234 226894 81854 238000
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 176600 81854 190338
rect 84954 230614 85574 238000
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 176600 85574 194058
rect 91794 237454 92414 238000
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 176600 92414 200898
rect 95514 205174 96134 238000
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 176600 96134 204618
rect 99234 208894 99854 238000
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 98315 177716 98381 177717
rect 98315 177652 98316 177716
rect 98380 177652 98381 177716
rect 98315 177651 98381 177652
rect 97027 177036 97093 177037
rect 97027 176972 97028 177036
rect 97092 176972 97093 177036
rect 97027 176971 97093 176972
rect 97030 175130 97090 176971
rect 96960 175070 97090 175130
rect 98318 175130 98378 177651
rect 99234 176600 99854 208338
rect 102954 212614 103574 238000
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 101995 176764 102061 176765
rect 101995 176700 101996 176764
rect 102060 176700 102061 176764
rect 101995 176699 102061 176700
rect 99419 176492 99485 176493
rect 99419 176428 99420 176492
rect 99484 176428 99485 176492
rect 99419 176427 99485 176428
rect 99422 175130 99482 176427
rect 100707 175404 100773 175405
rect 100707 175340 100708 175404
rect 100772 175340 100773 175404
rect 100707 175339 100773 175340
rect 98318 175070 98380 175130
rect 96960 174494 97020 175070
rect 98320 174494 98380 175070
rect 99408 175070 99482 175130
rect 100710 175130 100770 175339
rect 101998 175130 102058 176699
rect 102954 176600 103574 212058
rect 109794 219454 110414 238000
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 104571 177716 104637 177717
rect 104571 177652 104572 177716
rect 104636 177652 104637 177716
rect 104571 177651 104637 177652
rect 106963 177716 107029 177717
rect 106963 177652 106964 177716
rect 107028 177652 107029 177716
rect 106963 177651 107029 177652
rect 103283 176492 103349 176493
rect 103283 176428 103284 176492
rect 103348 176428 103349 176492
rect 103283 176427 103349 176428
rect 100710 175070 100828 175130
rect 99408 174494 99468 175070
rect 100768 174494 100828 175070
rect 101992 175070 102058 175130
rect 103286 175130 103346 176427
rect 104574 175130 104634 177651
rect 105675 176900 105741 176901
rect 105675 176836 105676 176900
rect 105740 176836 105741 176900
rect 105675 176835 105741 176836
rect 105678 175130 105738 176835
rect 103286 175070 103412 175130
rect 104574 175070 104636 175130
rect 101992 174494 102052 175070
rect 103352 174494 103412 175070
rect 104576 174494 104636 175070
rect 105664 175070 105738 175130
rect 106966 175130 107026 177651
rect 108067 176764 108133 176765
rect 108067 176700 108068 176764
rect 108132 176700 108133 176764
rect 108067 176699 108133 176700
rect 109539 176764 109605 176765
rect 109539 176700 109540 176764
rect 109604 176700 109605 176764
rect 109539 176699 109605 176700
rect 108070 175130 108130 176699
rect 109542 175130 109602 176699
rect 109794 176600 110414 182898
rect 113514 223174 114134 238000
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 110643 177716 110709 177717
rect 110643 177652 110644 177716
rect 110708 177652 110709 177716
rect 110643 177651 110709 177652
rect 106966 175070 107084 175130
rect 108070 175070 108172 175130
rect 105664 174494 105724 175070
rect 107024 174494 107084 175070
rect 108112 174494 108172 175070
rect 109472 175070 109602 175130
rect 110646 175130 110706 177651
rect 112115 177036 112181 177037
rect 112115 176972 112116 177036
rect 112180 176972 112181 177036
rect 112115 176971 112181 176972
rect 112118 175130 112178 176971
rect 113514 176600 114134 186618
rect 117234 226894 117854 238000
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 119294 219450 119354 240891
rect 124262 238509 124322 339355
rect 125734 238645 125794 343707
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 125731 238644 125797 238645
rect 125731 238580 125732 238644
rect 125796 238580 125797 238644
rect 125731 238579 125797 238580
rect 124259 238508 124325 238509
rect 124259 238444 124260 238508
rect 124324 238444 124325 238508
rect 124259 238443 124325 238444
rect 118926 219390 119354 219450
rect 120954 230614 121574 238000
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 118926 200701 118986 219390
rect 118923 200700 118989 200701
rect 118923 200636 118924 200700
rect 118988 200636 118989 200700
rect 118923 200635 118989 200636
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 114323 177716 114389 177717
rect 114323 177652 114324 177716
rect 114388 177652 114389 177716
rect 114323 177651 114389 177652
rect 115795 177716 115861 177717
rect 115795 177652 115796 177716
rect 115860 177652 115861 177716
rect 115795 177651 115861 177652
rect 116899 177716 116965 177717
rect 116899 177652 116900 177716
rect 116964 177652 116965 177716
rect 116899 177651 116965 177652
rect 113219 175540 113285 175541
rect 113219 175476 113220 175540
rect 113284 175476 113285 175540
rect 113219 175475 113285 175476
rect 113222 175130 113282 175475
rect 110646 175070 110756 175130
rect 109472 174494 109532 175070
rect 110696 174494 110756 175070
rect 112056 175070 112178 175130
rect 113144 175070 113282 175130
rect 114326 175130 114386 177651
rect 115798 175130 115858 177651
rect 114326 175070 114428 175130
rect 112056 174494 112116 175070
rect 113144 174494 113204 175070
rect 114368 174494 114428 175070
rect 115728 175070 115858 175130
rect 116902 175130 116962 177651
rect 117234 176600 117854 190338
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 119475 177716 119541 177717
rect 119475 177652 119476 177716
rect 119540 177652 119541 177716
rect 119475 177651 119541 177652
rect 120763 177716 120829 177717
rect 120763 177652 120764 177716
rect 120828 177652 120829 177716
rect 120763 177651 120829 177652
rect 118371 175404 118437 175405
rect 118371 175340 118372 175404
rect 118436 175340 118437 175404
rect 118371 175339 118437 175340
rect 118374 175130 118434 175339
rect 119478 175130 119538 177651
rect 120766 175130 120826 177651
rect 120954 176600 121574 194058
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 124443 177036 124509 177037
rect 124443 176972 124444 177036
rect 124508 176972 124509 177036
rect 124443 176971 124509 176972
rect 123155 176764 123221 176765
rect 123155 176700 123156 176764
rect 123220 176700 123221 176764
rect 123155 176699 123221 176700
rect 121867 175404 121933 175405
rect 121867 175340 121868 175404
rect 121932 175340 121933 175404
rect 121867 175339 121933 175340
rect 121870 175130 121930 175339
rect 123158 175130 123218 176699
rect 124446 175130 124506 176971
rect 125731 176764 125797 176765
rect 125731 176700 125732 176764
rect 125796 176700 125797 176764
rect 125731 176699 125797 176700
rect 125734 175130 125794 176699
rect 127794 176600 128414 200898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 129411 177716 129477 177717
rect 129411 177652 129412 177716
rect 129476 177652 129477 177716
rect 129411 177651 129477 177652
rect 130699 177716 130765 177717
rect 130699 177652 130700 177716
rect 130764 177652 130765 177716
rect 130699 177651 130765 177652
rect 128123 176492 128189 176493
rect 128123 176428 128124 176492
rect 128188 176428 128189 176492
rect 128123 176427 128189 176428
rect 127019 175540 127085 175541
rect 127019 175476 127020 175540
rect 127084 175476 127085 175540
rect 127019 175475 127085 175476
rect 127022 175130 127082 175475
rect 128126 175130 128186 176427
rect 116902 175070 117012 175130
rect 115728 174494 115788 175070
rect 116952 174494 117012 175070
rect 118312 175070 118434 175130
rect 119400 175070 119538 175130
rect 120760 175070 120826 175130
rect 121848 175070 121930 175130
rect 123072 175070 123218 175130
rect 124432 175070 124506 175130
rect 125656 175070 125794 175130
rect 127016 175070 127082 175130
rect 128104 175070 128186 175130
rect 129414 175130 129474 177651
rect 130702 175130 130762 177651
rect 131514 176600 132134 204618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 133091 176764 133157 176765
rect 133091 176700 133092 176764
rect 133156 176700 133157 176764
rect 133091 176699 133157 176700
rect 134379 176764 134445 176765
rect 134379 176700 134380 176764
rect 134444 176700 134445 176764
rect 134379 176699 134445 176700
rect 131987 175540 132053 175541
rect 131987 175476 131988 175540
rect 132052 175476 132053 175540
rect 131987 175475 132053 175476
rect 129414 175070 129524 175130
rect 118312 174494 118372 175070
rect 119400 174494 119460 175070
rect 120760 174494 120820 175070
rect 121848 174494 121908 175070
rect 123072 174494 123132 175070
rect 124432 174494 124492 175070
rect 125656 174494 125716 175070
rect 127016 174494 127076 175070
rect 128104 174494 128164 175070
rect 129464 174494 129524 175070
rect 130688 175070 130762 175130
rect 131990 175130 132050 175475
rect 133094 175130 133154 176699
rect 134382 175130 134442 176699
rect 135234 176600 135854 208338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 136035 176764 136101 176765
rect 136035 176700 136036 176764
rect 136100 176700 136101 176764
rect 136035 176699 136101 176700
rect 136038 175130 136098 176699
rect 138954 176600 139574 212058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 176600 146414 182898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 148179 176764 148245 176765
rect 148179 176700 148180 176764
rect 148244 176700 148245 176764
rect 148179 176699 148245 176700
rect 131990 175070 132108 175130
rect 133094 175070 133196 175130
rect 130688 174494 130748 175070
rect 132048 174494 132108 175070
rect 133136 174494 133196 175070
rect 134360 175070 134442 175130
rect 135720 175070 136098 175130
rect 148182 175130 148242 176699
rect 149514 176600 150134 186618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 176600 153854 190338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 176600 157574 194058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 176600 164414 200898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 170259 381308 170325 381309
rect 170259 381244 170260 381308
rect 170324 381244 170325 381308
rect 170259 381243 170325 381244
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 166211 179484 166277 179485
rect 166211 179420 166212 179484
rect 166276 179420 166277 179484
rect 166211 179419 166277 179420
rect 158851 175540 158917 175541
rect 158851 175476 158852 175540
rect 158916 175476 158917 175540
rect 158851 175475 158917 175476
rect 158854 175130 158914 175475
rect 148182 175070 148292 175130
rect 134360 174494 134420 175070
rect 135720 174494 135780 175070
rect 148232 174494 148292 175070
rect 158840 175070 158914 175130
rect 158840 174494 158900 175070
rect 69072 165454 69420 165486
rect 69072 165218 69128 165454
rect 69364 165218 69420 165454
rect 69072 165134 69420 165218
rect 69072 164898 69128 165134
rect 69364 164898 69420 165134
rect 69072 164866 69420 164898
rect 164136 165454 164484 165486
rect 164136 165218 164192 165454
rect 164428 165218 164484 165454
rect 164136 165134 164484 165218
rect 164136 164898 164192 165134
rect 164428 164898 164484 165134
rect 164136 164866 164484 164898
rect 166214 154597 166274 179419
rect 166395 175404 166461 175405
rect 166395 175340 166396 175404
rect 166460 175340 166461 175404
rect 166395 175339 166461 175340
rect 166398 163165 166458 175339
rect 167514 169174 168134 204618
rect 168235 176900 168301 176901
rect 168235 176836 168236 176900
rect 168300 176836 168301 176900
rect 168235 176835 168301 176836
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 166395 163164 166461 163165
rect 166395 163100 166396 163164
rect 166460 163100 166461 163164
rect 166395 163099 166461 163100
rect 166211 154596 166277 154597
rect 166211 154532 166212 154596
rect 166276 154532 166277 154596
rect 166211 154531 166277 154532
rect 69752 147454 70100 147486
rect 69752 147218 69808 147454
rect 70044 147218 70100 147454
rect 69752 147134 70100 147218
rect 69752 146898 69808 147134
rect 70044 146898 70100 147134
rect 69752 146866 70100 146898
rect 163456 147454 163804 147486
rect 163456 147218 163512 147454
rect 163748 147218 163804 147454
rect 163456 147134 163804 147218
rect 163456 146898 163512 147134
rect 163748 146898 163804 147134
rect 163456 146866 163804 146898
rect 166395 134196 166461 134197
rect 166395 134132 166396 134196
rect 166460 134132 166461 134196
rect 166395 134131 166461 134132
rect 166211 130116 166277 130117
rect 166211 130052 166212 130116
rect 166276 130052 166277 130116
rect 166211 130051 166277 130052
rect 69072 129454 69420 129486
rect 69072 129218 69128 129454
rect 69364 129218 69420 129454
rect 69072 129134 69420 129218
rect 69072 128898 69128 129134
rect 69364 128898 69420 129134
rect 69072 128866 69420 128898
rect 164136 129454 164484 129486
rect 164136 129218 164192 129454
rect 164428 129218 164484 129454
rect 164136 129134 164484 129218
rect 164136 128898 164192 129134
rect 164428 128898 164484 129134
rect 164136 128866 164484 128898
rect 69752 111454 70100 111486
rect 69752 111218 69808 111454
rect 70044 111218 70100 111454
rect 69752 111134 70100 111218
rect 69752 110898 69808 111134
rect 70044 110898 70100 111134
rect 69752 110866 70100 110898
rect 163456 111454 163804 111486
rect 163456 111218 163512 111454
rect 163748 111218 163804 111454
rect 163456 111134 163804 111218
rect 163456 110898 163512 111134
rect 163748 110898 163804 111134
rect 163456 110866 163804 110898
rect 74656 94890 74716 95200
rect 84312 94890 84372 95200
rect 85536 94890 85596 95200
rect 86624 94890 86684 95200
rect 87984 94890 88044 95200
rect 88936 94890 88996 95200
rect 74656 94830 74826 94890
rect 84312 94830 84394 94890
rect 85536 94830 85682 94890
rect 86624 94830 86786 94890
rect 87984 94830 88074 94890
rect 66954 68614 67574 93100
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 66115 13156 66181 13157
rect 66115 13092 66116 13156
rect 66180 13092 66181 13156
rect 66115 13091 66181 13092
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 75454 74414 93100
rect 74766 92445 74826 94830
rect 74763 92444 74829 92445
rect 74763 92380 74764 92444
rect 74828 92380 74829 92444
rect 74763 92379 74829 92380
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 79174 78134 93100
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 82894 81854 93100
rect 84334 91221 84394 94830
rect 85622 93669 85682 94830
rect 85619 93668 85685 93669
rect 85619 93604 85620 93668
rect 85684 93604 85685 93668
rect 85619 93603 85685 93604
rect 84331 91220 84397 91221
rect 84331 91156 84332 91220
rect 84396 91156 84397 91220
rect 84331 91155 84397 91156
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 86614 85574 93100
rect 86726 91221 86786 94830
rect 88014 91221 88074 94830
rect 88934 94830 88996 94890
rect 90160 94890 90220 95200
rect 91384 94890 91444 95200
rect 90160 94830 90282 94890
rect 88934 92445 88994 94830
rect 88931 92444 88997 92445
rect 88931 92380 88932 92444
rect 88996 92380 88997 92444
rect 88931 92379 88997 92380
rect 90222 91221 90282 94830
rect 91326 94830 91444 94890
rect 92472 94890 92532 95200
rect 93832 94890 93892 95200
rect 94920 94890 94980 95200
rect 96008 94890 96068 95200
rect 96688 94890 96748 95200
rect 92472 94830 92674 94890
rect 93832 94830 93962 94890
rect 94920 94830 95066 94890
rect 96008 94830 96354 94890
rect 91326 91221 91386 94830
rect 86723 91220 86789 91221
rect 86723 91156 86724 91220
rect 86788 91156 86789 91220
rect 86723 91155 86789 91156
rect 88011 91220 88077 91221
rect 88011 91156 88012 91220
rect 88076 91156 88077 91220
rect 88011 91155 88077 91156
rect 90219 91220 90285 91221
rect 90219 91156 90220 91220
rect 90284 91156 90285 91220
rect 90219 91155 90285 91156
rect 91323 91220 91389 91221
rect 91323 91156 91324 91220
rect 91388 91156 91389 91220
rect 91323 91155 91389 91156
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 93100
rect 92614 91221 92674 94830
rect 93902 91221 93962 94830
rect 95006 92445 95066 94830
rect 95003 92444 95069 92445
rect 95003 92380 95004 92444
rect 95068 92380 95069 92444
rect 95003 92379 95069 92380
rect 92611 91220 92677 91221
rect 92611 91156 92612 91220
rect 92676 91156 92677 91220
rect 92611 91155 92677 91156
rect 93899 91220 93965 91221
rect 93899 91156 93900 91220
rect 93964 91156 93965 91220
rect 93899 91155 93965 91156
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 61174 96134 93100
rect 96294 91221 96354 94830
rect 96662 94830 96748 94890
rect 97096 94890 97156 95200
rect 98048 94890 98108 95200
rect 98456 94890 98516 95200
rect 99136 94890 99196 95200
rect 97096 94830 97274 94890
rect 98048 94830 98194 94890
rect 98456 94830 98562 94890
rect 96662 91221 96722 94830
rect 97214 91221 97274 94830
rect 98134 91221 98194 94830
rect 98502 91357 98562 94830
rect 99054 94830 99196 94890
rect 99544 94890 99604 95200
rect 100632 94890 100692 95200
rect 99544 94830 100034 94890
rect 98499 91356 98565 91357
rect 98499 91292 98500 91356
rect 98564 91292 98565 91356
rect 98499 91291 98565 91292
rect 99054 91221 99114 94830
rect 96291 91220 96357 91221
rect 96291 91156 96292 91220
rect 96356 91156 96357 91220
rect 96291 91155 96357 91156
rect 96659 91220 96725 91221
rect 96659 91156 96660 91220
rect 96724 91156 96725 91220
rect 96659 91155 96725 91156
rect 97211 91220 97277 91221
rect 97211 91156 97212 91220
rect 97276 91156 97277 91220
rect 97211 91155 97277 91156
rect 98131 91220 98197 91221
rect 98131 91156 98132 91220
rect 98196 91156 98197 91220
rect 98131 91155 98197 91156
rect 99051 91220 99117 91221
rect 99051 91156 99052 91220
rect 99116 91156 99117 91220
rect 99051 91155 99117 91156
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 64894 99854 93100
rect 99974 91221 100034 94830
rect 100526 94830 100692 94890
rect 100768 94890 100828 95200
rect 101856 94890 101916 95200
rect 100768 94830 100954 94890
rect 100526 91221 100586 94830
rect 100894 91357 100954 94830
rect 101814 94830 101916 94890
rect 101992 94890 102052 95200
rect 102944 94890 103004 95200
rect 101992 94830 102058 94890
rect 101814 92445 101874 94830
rect 101811 92444 101877 92445
rect 101811 92380 101812 92444
rect 101876 92380 101877 92444
rect 101811 92379 101877 92380
rect 100891 91356 100957 91357
rect 100891 91292 100892 91356
rect 100956 91292 100957 91356
rect 100891 91291 100957 91292
rect 101998 91221 102058 94830
rect 102918 94830 103004 94890
rect 103216 94890 103276 95200
rect 104304 94890 104364 95200
rect 103216 94830 103346 94890
rect 102918 93870 102978 94830
rect 102734 93810 102978 93870
rect 102734 91221 102794 93810
rect 103286 93261 103346 94830
rect 104206 94830 104364 94890
rect 104440 94890 104500 95200
rect 105392 94890 105452 95200
rect 105664 94890 105724 95200
rect 104440 94830 104634 94890
rect 105392 94830 105554 94890
rect 105664 94830 105738 94890
rect 103283 93260 103349 93261
rect 103283 93196 103284 93260
rect 103348 93196 103349 93260
rect 103283 93195 103349 93196
rect 99971 91220 100037 91221
rect 99971 91156 99972 91220
rect 100036 91156 100037 91220
rect 99971 91155 100037 91156
rect 100523 91220 100589 91221
rect 100523 91156 100524 91220
rect 100588 91156 100589 91220
rect 100523 91155 100589 91156
rect 101995 91220 102061 91221
rect 101995 91156 101996 91220
rect 102060 91156 102061 91220
rect 101995 91155 102061 91156
rect 102731 91220 102797 91221
rect 102731 91156 102732 91220
rect 102796 91156 102797 91220
rect 102731 91155 102797 91156
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 68614 103574 93100
rect 104206 91357 104266 94830
rect 104203 91356 104269 91357
rect 104203 91292 104204 91356
rect 104268 91292 104269 91356
rect 104203 91291 104269 91292
rect 104574 91221 104634 94830
rect 105494 92445 105554 94830
rect 105491 92444 105557 92445
rect 105491 92380 105492 92444
rect 105556 92380 105557 92444
rect 105491 92379 105557 92380
rect 105678 91765 105738 94830
rect 106227 94756 106293 94757
rect 106227 94692 106228 94756
rect 106292 94692 106293 94756
rect 106227 94691 106293 94692
rect 106230 92445 106290 94691
rect 106480 94210 106540 95200
rect 106616 94757 106676 95200
rect 107704 94890 107764 95200
rect 108112 94890 108172 95200
rect 107702 94830 107764 94890
rect 108070 94830 108172 94890
rect 109064 94890 109124 95200
rect 109472 94890 109532 95200
rect 110152 94890 110212 95200
rect 110696 94890 110756 95200
rect 111240 94890 111300 95200
rect 109064 94830 109234 94890
rect 109472 94830 109602 94890
rect 110152 94830 110338 94890
rect 106613 94756 106679 94757
rect 106613 94692 106614 94756
rect 106678 94692 106679 94756
rect 106613 94691 106679 94692
rect 106480 94150 106658 94210
rect 106227 92444 106293 92445
rect 106227 92380 106228 92444
rect 106292 92380 106293 92444
rect 106227 92379 106293 92380
rect 105675 91764 105741 91765
rect 105675 91700 105676 91764
rect 105740 91700 105741 91764
rect 105675 91699 105741 91700
rect 106598 91221 106658 94150
rect 107702 91221 107762 94830
rect 108070 91357 108130 94830
rect 108067 91356 108133 91357
rect 108067 91292 108068 91356
rect 108132 91292 108133 91356
rect 108067 91291 108133 91292
rect 109174 91221 109234 94830
rect 109542 91357 109602 94830
rect 110278 93261 110338 94830
rect 110646 94830 110756 94890
rect 111198 94830 111300 94890
rect 111920 94890 111980 95200
rect 112328 94890 112388 95200
rect 111920 94830 111994 94890
rect 110275 93260 110341 93261
rect 110275 93196 110276 93260
rect 110340 93196 110341 93260
rect 110275 93195 110341 93196
rect 109539 91356 109605 91357
rect 109539 91292 109540 91356
rect 109604 91292 109605 91356
rect 109539 91291 109605 91292
rect 104571 91220 104637 91221
rect 104571 91156 104572 91220
rect 104636 91156 104637 91220
rect 104571 91155 104637 91156
rect 106595 91220 106661 91221
rect 106595 91156 106596 91220
rect 106660 91156 106661 91220
rect 106595 91155 106661 91156
rect 107699 91220 107765 91221
rect 107699 91156 107700 91220
rect 107764 91156 107765 91220
rect 107699 91155 107765 91156
rect 109171 91220 109237 91221
rect 109171 91156 109172 91220
rect 109236 91156 109237 91220
rect 109171 91155 109237 91156
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 75454 110414 93100
rect 110646 91221 110706 94830
rect 111198 91221 111258 94830
rect 111934 93941 111994 94830
rect 112302 94830 112388 94890
rect 113144 94890 113204 95200
rect 113688 94890 113748 95200
rect 114368 94890 114428 95200
rect 113144 94830 113282 94890
rect 113688 94830 113834 94890
rect 111931 93940 111997 93941
rect 111931 93876 111932 93940
rect 111996 93876 111997 93940
rect 111931 93875 111997 93876
rect 112302 91221 112362 94830
rect 113222 91221 113282 94830
rect 113774 93261 113834 94830
rect 114326 94830 114428 94890
rect 114776 94890 114836 95200
rect 115456 94890 115516 95200
rect 115864 94890 115924 95200
rect 114776 94830 114938 94890
rect 113771 93260 113837 93261
rect 113771 93196 113772 93260
rect 113836 93196 113837 93260
rect 113771 93195 113837 93196
rect 110643 91220 110709 91221
rect 110643 91156 110644 91220
rect 110708 91156 110709 91220
rect 110643 91155 110709 91156
rect 111195 91220 111261 91221
rect 111195 91156 111196 91220
rect 111260 91156 111261 91220
rect 111195 91155 111261 91156
rect 112299 91220 112365 91221
rect 112299 91156 112300 91220
rect 112364 91156 112365 91220
rect 112299 91155 112365 91156
rect 113219 91220 113285 91221
rect 113219 91156 113220 91220
rect 113284 91156 113285 91220
rect 113219 91155 113285 91156
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 79174 114134 93100
rect 114326 92309 114386 94830
rect 114323 92308 114389 92309
rect 114323 92244 114324 92308
rect 114388 92244 114389 92308
rect 114323 92243 114389 92244
rect 114878 91765 114938 94830
rect 115430 94830 115516 94890
rect 115798 94830 115924 94890
rect 116680 94890 116740 95200
rect 117088 94890 117148 95200
rect 116680 94830 116778 94890
rect 115430 93669 115490 94830
rect 115427 93668 115493 93669
rect 115427 93604 115428 93668
rect 115492 93604 115493 93668
rect 115427 93603 115493 93604
rect 114875 91764 114941 91765
rect 114875 91700 114876 91764
rect 114940 91700 114941 91764
rect 114875 91699 114941 91700
rect 115798 91221 115858 94830
rect 116718 92445 116778 94830
rect 117086 94830 117148 94890
rect 117904 94890 117964 95200
rect 118176 94890 118236 95200
rect 119400 94890 119460 95200
rect 117904 94830 118066 94890
rect 118176 94830 118250 94890
rect 116715 92444 116781 92445
rect 116715 92380 116716 92444
rect 116780 92380 116781 92444
rect 116715 92379 116781 92380
rect 117086 91221 117146 94830
rect 115795 91220 115861 91221
rect 115795 91156 115796 91220
rect 115860 91156 115861 91220
rect 115795 91155 115861 91156
rect 117083 91220 117149 91221
rect 117083 91156 117084 91220
rect 117148 91156 117149 91220
rect 117083 91155 117149 91156
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 82894 117854 93100
rect 118006 91221 118066 94830
rect 118190 91357 118250 94830
rect 119294 94830 119460 94890
rect 119536 94890 119596 95200
rect 120216 94890 120276 95200
rect 120624 94890 120684 95200
rect 121712 94890 121772 95200
rect 119536 94830 119722 94890
rect 119294 91357 119354 94830
rect 118187 91356 118253 91357
rect 118187 91292 118188 91356
rect 118252 91292 118253 91356
rect 118187 91291 118253 91292
rect 119291 91356 119357 91357
rect 119291 91292 119292 91356
rect 119356 91292 119357 91356
rect 119291 91291 119357 91292
rect 119662 91221 119722 94830
rect 120214 94830 120276 94890
rect 120582 94830 120684 94890
rect 121686 94830 121772 94890
rect 121984 94890 122044 95200
rect 122800 94890 122860 95200
rect 123208 94890 123268 95200
rect 121984 94830 122114 94890
rect 122800 94830 123034 94890
rect 120214 91221 120274 94830
rect 120582 93669 120642 94830
rect 120579 93668 120645 93669
rect 120579 93604 120580 93668
rect 120644 93604 120645 93668
rect 120579 93603 120645 93604
rect 118003 91220 118069 91221
rect 118003 91156 118004 91220
rect 118068 91156 118069 91220
rect 118003 91155 118069 91156
rect 119659 91220 119725 91221
rect 119659 91156 119660 91220
rect 119724 91156 119725 91220
rect 119659 91155 119725 91156
rect 120211 91220 120277 91221
rect 120211 91156 120212 91220
rect 120276 91156 120277 91220
rect 120211 91155 120277 91156
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 86614 121574 93100
rect 121686 91357 121746 94830
rect 121683 91356 121749 91357
rect 121683 91292 121684 91356
rect 121748 91292 121749 91356
rect 121683 91291 121749 91292
rect 122054 91221 122114 94830
rect 122974 93870 123034 94830
rect 122606 93810 123034 93870
rect 123158 94830 123268 94890
rect 124024 94890 124084 95200
rect 124432 94890 124492 95200
rect 125384 94890 125444 95200
rect 124024 94830 124138 94890
rect 124432 94830 124506 94890
rect 122606 91490 122666 93810
rect 122787 91492 122853 91493
rect 122787 91490 122788 91492
rect 122606 91430 122788 91490
rect 122787 91428 122788 91430
rect 122852 91428 122853 91492
rect 122787 91427 122853 91428
rect 123158 91221 123218 94830
rect 124078 92445 124138 94830
rect 124075 92444 124141 92445
rect 124075 92380 124076 92444
rect 124140 92380 124141 92444
rect 124075 92379 124141 92380
rect 124446 91629 124506 94830
rect 125366 94830 125444 94890
rect 125656 94890 125716 95200
rect 126472 94890 126532 95200
rect 125656 94830 125794 94890
rect 124443 91628 124509 91629
rect 124443 91564 124444 91628
rect 124508 91564 124509 91628
rect 124443 91563 124509 91564
rect 125366 91221 125426 94830
rect 125734 92445 125794 94830
rect 126470 94830 126532 94890
rect 126608 94890 126668 95200
rect 128104 94890 128164 95200
rect 126608 94830 126714 94890
rect 128104 94830 128186 94890
rect 125731 92444 125797 92445
rect 125731 92380 125732 92444
rect 125796 92380 125797 92444
rect 125731 92379 125797 92380
rect 126470 91629 126530 94830
rect 126654 92037 126714 94830
rect 128126 93261 128186 94830
rect 129328 94757 129388 95200
rect 130688 94890 130748 95200
rect 131912 94890 131972 95200
rect 133136 94890 133196 95200
rect 130688 94830 130762 94890
rect 131912 94830 132418 94890
rect 129325 94756 129391 94757
rect 129325 94692 129326 94756
rect 129390 94692 129391 94756
rect 129325 94691 129391 94692
rect 128123 93260 128189 93261
rect 128123 93196 128124 93260
rect 128188 93196 128189 93260
rect 128123 93195 128189 93196
rect 126651 92036 126717 92037
rect 126651 91972 126652 92036
rect 126716 91972 126717 92036
rect 126651 91971 126717 91972
rect 126467 91628 126533 91629
rect 126467 91564 126468 91628
rect 126532 91564 126533 91628
rect 126467 91563 126533 91564
rect 122051 91220 122117 91221
rect 122051 91156 122052 91220
rect 122116 91156 122117 91220
rect 122051 91155 122117 91156
rect 123155 91220 123221 91221
rect 123155 91156 123156 91220
rect 123220 91156 123221 91220
rect 123155 91155 123221 91156
rect 125363 91220 125429 91221
rect 125363 91156 125364 91220
rect 125428 91156 125429 91220
rect 125363 91155 125429 91156
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 93100
rect 130702 91221 130762 94830
rect 130699 91220 130765 91221
rect 130699 91156 130700 91220
rect 130764 91156 130765 91220
rect 130699 91155 130765 91156
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 61174 132134 93100
rect 132358 91221 132418 94830
rect 133094 94830 133196 94890
rect 134360 94890 134420 95200
rect 135584 94890 135644 95200
rect 151496 94890 151556 95200
rect 134360 94830 134442 94890
rect 135584 94830 135730 94890
rect 133094 91221 133154 94830
rect 134382 92445 134442 94830
rect 135670 93669 135730 94830
rect 151494 94830 151556 94890
rect 135667 93668 135733 93669
rect 135667 93604 135668 93668
rect 135732 93604 135733 93668
rect 135667 93603 135733 93604
rect 134379 92444 134445 92445
rect 134379 92380 134380 92444
rect 134444 92380 134445 92444
rect 134379 92379 134445 92380
rect 132355 91220 132421 91221
rect 132355 91156 132356 91220
rect 132420 91156 132421 91220
rect 132355 91155 132421 91156
rect 133091 91220 133157 91221
rect 133091 91156 133092 91220
rect 133156 91156 133157 91220
rect 133091 91155 133157 91156
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 64894 135854 93100
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 68614 139574 93100
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 75454 146414 93100
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 79174 150134 93100
rect 151494 91221 151554 94830
rect 151632 94210 151692 95200
rect 151768 94757 151828 95200
rect 151904 94890 151964 95200
rect 151904 94830 152106 94890
rect 151765 94756 151831 94757
rect 151765 94692 151766 94756
rect 151830 94692 151831 94756
rect 151765 94691 151831 94692
rect 151632 94150 151738 94210
rect 151678 93669 151738 94150
rect 151675 93668 151741 93669
rect 151675 93604 151676 93668
rect 151740 93604 151741 93668
rect 151675 93603 151741 93604
rect 152046 92445 152106 94830
rect 152043 92444 152109 92445
rect 152043 92380 152044 92444
rect 152108 92380 152109 92444
rect 152043 92379 152109 92380
rect 151491 91220 151557 91221
rect 151491 91156 151492 91220
rect 151556 91156 151557 91220
rect 151491 91155 151557 91156
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 82894 153854 93100
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 86614 157574 93100
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 93100
rect 166214 84149 166274 130051
rect 166398 88229 166458 134131
rect 167514 133174 168134 168618
rect 168238 158813 168298 176835
rect 168235 158812 168301 158813
rect 168235 158748 168236 158812
rect 168300 158748 168301 158812
rect 168235 158747 168301 158748
rect 169155 135284 169221 135285
rect 169155 135220 169156 135284
rect 169220 135220 169221 135284
rect 169155 135219 169221 135220
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 168971 128620 169037 128621
rect 168971 128556 168972 128620
rect 169036 128556 169037 128620
rect 168971 128555 169037 128556
rect 168235 127124 168301 127125
rect 168235 127060 168236 127124
rect 168300 127060 168301 127124
rect 168235 127059 168301 127060
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 166395 88228 166461 88229
rect 166395 88164 166396 88228
rect 166460 88164 166461 88228
rect 166395 88163 166461 88164
rect 166211 84148 166277 84149
rect 166211 84084 166212 84148
rect 166276 84084 166277 84148
rect 166211 84083 166277 84084
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 61174 168134 96618
rect 168238 91085 168298 127059
rect 168235 91084 168301 91085
rect 168235 91020 168236 91084
rect 168300 91020 168301 91084
rect 168235 91019 168301 91020
rect 168974 80069 169034 128555
rect 169158 93941 169218 135219
rect 170262 115157 170322 381243
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 170443 138140 170509 138141
rect 170443 138076 170444 138140
rect 170508 138076 170509 138140
rect 170443 138075 170509 138076
rect 170259 115156 170325 115157
rect 170259 115092 170260 115156
rect 170324 115092 170325 115156
rect 170259 115091 170325 115092
rect 170259 99516 170325 99517
rect 170259 99452 170260 99516
rect 170324 99452 170325 99516
rect 170259 99451 170325 99452
rect 169155 93940 169221 93941
rect 169155 93876 169156 93940
rect 169220 93876 169221 93940
rect 169155 93875 169221 93876
rect 170262 86869 170322 99451
rect 170259 86868 170325 86869
rect 170259 86804 170260 86868
rect 170324 86804 170325 86868
rect 170259 86803 170325 86804
rect 170446 84013 170506 138075
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 177251 387836 177317 387837
rect 177251 387772 177252 387836
rect 177316 387772 177317 387836
rect 177251 387771 177317 387772
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 173019 105228 173085 105229
rect 173019 105164 173020 105228
rect 173084 105164 173085 105228
rect 173019 105163 173085 105164
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 170443 84012 170509 84013
rect 170443 83948 170444 84012
rect 170508 83948 170509 84012
rect 170443 83947 170509 83948
rect 168971 80068 169037 80069
rect 168971 80004 168972 80068
rect 169036 80004 169037 80068
rect 168971 80003 169037 80004
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 64894 171854 100338
rect 173022 94893 173082 105163
rect 174954 104614 175574 140058
rect 177254 106861 177314 387771
rect 178539 373692 178605 373693
rect 178539 373628 178540 373692
rect 178604 373628 178605 373692
rect 178539 373627 178605 373628
rect 177251 106860 177317 106861
rect 177251 106796 177252 106860
rect 177316 106796 177317 106860
rect 177251 106795 177317 106796
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 173019 94892 173085 94893
rect 173019 94828 173020 94892
rect 173084 94828 173085 94892
rect 173019 94827 173085 94828
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 68614 175574 104058
rect 178542 80749 178602 373627
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 178539 80748 178605 80749
rect 178539 80684 178540 80748
rect 178604 80684 178605 80748
rect 178539 80683 178605 80684
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 277174 204134 312618
rect 203514 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 204134 277174
rect 203514 276854 204134 276938
rect 203514 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 204134 276854
rect 203514 241174 204134 276618
rect 203514 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 204134 241174
rect 203514 240854 204134 240938
rect 203514 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 204134 240854
rect 203514 205174 204134 240618
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 280894 207854 316338
rect 207234 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 207854 280894
rect 207234 280574 207854 280658
rect 207234 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 207854 280574
rect 207234 244894 207854 280338
rect 207234 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 207854 244894
rect 207234 244574 207854 244658
rect 207234 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 207854 244574
rect 207234 208894 207854 244338
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 284614 211574 320058
rect 210954 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 211574 284614
rect 210954 284294 211574 284378
rect 210954 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 211574 284294
rect 210954 248614 211574 284058
rect 210954 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 211574 248614
rect 210954 248294 211574 248378
rect 210954 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 211574 248294
rect 210954 212614 211574 248058
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 178000 218414 182898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 223174 222134 258618
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 178000 222134 186618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 262894 225854 298338
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 226894 225854 262338
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 178000 225854 190338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 266614 229574 302058
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228954 230614 229574 266058
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 178000 229574 194058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 178000 236414 200898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385174 240134 420618
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 349174 240134 384618
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 239514 313174 240134 348618
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 239514 277174 240134 312618
rect 239514 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 240134 277174
rect 239514 276854 240134 276938
rect 239514 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 240134 276854
rect 239514 241174 240134 276618
rect 239514 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 240134 241174
rect 239514 240854 240134 240938
rect 239514 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 240134 240854
rect 239514 205174 240134 240618
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 239514 178000 240134 204618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 352894 243854 388338
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 243234 316894 243854 352338
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 243234 280894 243854 316338
rect 243234 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 243854 280894
rect 243234 280574 243854 280658
rect 243234 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 243854 280574
rect 243234 244894 243854 280338
rect 243234 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 243854 244894
rect 243234 244574 243854 244658
rect 243234 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 243854 244574
rect 243234 208894 243854 244338
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 243234 178000 243854 208338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 356614 247574 392058
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 246954 320614 247574 356058
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 246954 284614 247574 320058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 252507 295492 252573 295493
rect 252507 295428 252508 295492
rect 252572 295428 252573 295492
rect 252507 295427 252573 295428
rect 246954 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 247574 284614
rect 246954 284294 247574 284378
rect 246954 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 247574 284294
rect 246954 248614 247574 284058
rect 246954 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 247574 248614
rect 246954 248294 247574 248378
rect 246954 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 247574 248294
rect 246954 212614 247574 248058
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 246954 178000 247574 212058
rect 249195 177580 249261 177581
rect 249195 177516 249196 177580
rect 249260 177516 249261 177580
rect 249195 177515 249261 177516
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 140614 211574 176058
rect 249198 174725 249258 177515
rect 249379 177444 249445 177445
rect 249379 177380 249380 177444
rect 249444 177380 249445 177444
rect 249379 177379 249445 177380
rect 249195 174724 249261 174725
rect 249195 174660 249196 174724
rect 249260 174660 249261 174724
rect 249195 174659 249261 174660
rect 249382 173365 249442 177379
rect 249379 173364 249445 173365
rect 249379 173300 249380 173364
rect 249444 173300 249445 173364
rect 249379 173299 249445 173300
rect 227874 165454 228194 165486
rect 227874 165218 227916 165454
rect 228152 165218 228194 165454
rect 227874 165134 228194 165218
rect 227874 164898 227916 165134
rect 228152 164898 228194 165134
rect 227874 164866 228194 164898
rect 237805 165454 238125 165486
rect 237805 165218 237847 165454
rect 238083 165218 238125 165454
rect 237805 165134 238125 165218
rect 237805 164898 237847 165134
rect 238083 164898 238125 165134
rect 237805 164866 238125 164898
rect 222910 147454 223230 147486
rect 222910 147218 222952 147454
rect 223188 147218 223230 147454
rect 222910 147134 223230 147218
rect 222910 146898 222952 147134
rect 223188 146898 223230 147134
rect 222910 146866 223230 146898
rect 232840 147454 233160 147486
rect 232840 147218 232882 147454
rect 233118 147218 233160 147454
rect 232840 147134 233160 147218
rect 232840 146898 232882 147134
rect 233118 146898 233160 147134
rect 232840 146866 233160 146898
rect 242771 147454 243091 147486
rect 242771 147218 242813 147454
rect 243049 147218 243091 147454
rect 242771 147134 243091 147218
rect 242771 146898 242813 147134
rect 243049 146898 243091 147134
rect 242771 146866 243091 146898
rect 251771 142764 251837 142765
rect 251771 142700 251772 142764
rect 251836 142700 251837 142764
rect 251771 142699 251837 142700
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 227874 129454 228194 129486
rect 227874 129218 227916 129454
rect 228152 129218 228194 129454
rect 227874 129134 228194 129218
rect 227874 128898 227916 129134
rect 228152 128898 228194 129134
rect 227874 128866 228194 128898
rect 237805 129454 238125 129486
rect 237805 129218 237847 129454
rect 238083 129218 238125 129454
rect 237805 129134 238125 129218
rect 237805 128898 237847 129134
rect 238083 128898 238125 129134
rect 237805 128866 238125 128898
rect 222910 111454 223230 111486
rect 222910 111218 222952 111454
rect 223188 111218 223230 111454
rect 222910 111134 223230 111218
rect 222910 110898 222952 111134
rect 223188 110898 223230 111134
rect 222910 110866 223230 110898
rect 232840 111454 233160 111486
rect 232840 111218 232882 111454
rect 233118 111218 233160 111454
rect 232840 111134 233160 111218
rect 232840 110898 232882 111134
rect 233118 110898 233160 111134
rect 232840 110866 233160 110898
rect 242771 111454 243091 111486
rect 242771 111218 242813 111454
rect 243049 111218 243091 111454
rect 242771 111134 243091 111218
rect 242771 110898 242813 111134
rect 243049 110898 243091 111134
rect 242771 110866 243091 110898
rect 214603 105092 214669 105093
rect 214603 105028 214604 105092
rect 214668 105028 214669 105092
rect 214603 105027 214669 105028
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 214419 97068 214485 97069
rect 214419 97004 214420 97068
rect 214484 97004 214485 97068
rect 214419 97003 214485 97004
rect 214422 81429 214482 97003
rect 214606 93805 214666 105027
rect 251774 104685 251834 142699
rect 252510 138005 252570 295427
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 259499 379132 259565 379133
rect 259499 379068 259500 379132
rect 259564 379068 259565 379132
rect 259499 379067 259565 379068
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 295174 258134 330618
rect 258395 301476 258461 301477
rect 258395 301412 258396 301476
rect 258460 301412 258461 301476
rect 258395 301411 258461 301412
rect 258398 296730 258458 301411
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 255267 274684 255333 274685
rect 255267 274620 255268 274684
rect 255332 274620 255333 274684
rect 255267 274619 255333 274620
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 255270 152149 255330 274619
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 223174 258134 258618
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 256739 185604 256805 185605
rect 256739 185540 256740 185604
rect 256804 185540 256805 185604
rect 256739 185539 256805 185540
rect 255267 152148 255333 152149
rect 255267 152084 255268 152148
rect 255332 152084 255333 152148
rect 255267 152083 255333 152084
rect 256742 147525 256802 185539
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 256739 147524 256805 147525
rect 256739 147460 256740 147524
rect 256804 147460 256805 147524
rect 256739 147459 256805 147460
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 252507 138004 252573 138005
rect 252507 137940 252508 138004
rect 252572 137940 252573 138004
rect 252507 137939 252573 137940
rect 253059 134196 253125 134197
rect 253059 134132 253060 134196
rect 253124 134132 253125 134196
rect 253059 134131 253125 134132
rect 251771 104684 251837 104685
rect 251771 104620 251772 104684
rect 251836 104620 251837 104684
rect 251771 104619 251837 104620
rect 214603 93804 214669 93805
rect 214603 93740 214604 93804
rect 214668 93740 214669 93804
rect 214603 93739 214669 93740
rect 214419 81428 214485 81429
rect 214419 81364 214420 81428
rect 214484 81364 214485 81428
rect 214419 81363 214485 81364
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 75454 218414 94000
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 79174 222134 94000
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 82894 225854 94000
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 86614 229574 94000
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 93454 236414 94000
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 61174 240134 94000
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 64894 243854 94000
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 68614 247574 94000
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253062 19957 253122 134131
rect 253794 111454 254414 146898
rect 254531 141540 254597 141541
rect 254531 141476 254532 141540
rect 254596 141476 254597 141540
rect 254531 141475 254597 141476
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 254534 101829 254594 141475
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 254531 101828 254597 101829
rect 254531 101764 254532 101828
rect 254596 101764 254597 101828
rect 254531 101763 254597 101764
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253059 19956 253125 19957
rect 253059 19892 253060 19956
rect 253124 19892 253125 19956
rect 253059 19891 253125 19892
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 258214 296670 258458 296730
rect 258214 16590 258274 296670
rect 258395 218652 258461 218653
rect 258395 218588 258396 218652
rect 258460 218588 258461 218652
rect 258395 218587 258461 218588
rect 258398 159357 258458 218587
rect 258395 159356 258461 159357
rect 258395 159292 258396 159356
rect 258460 159292 258461 159356
rect 258395 159291 258461 159292
rect 258214 16530 258458 16590
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 258398 3501 258458 16530
rect 259502 3501 259562 379067
rect 261234 370894 261854 406338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 262811 381172 262877 381173
rect 262811 381108 262812 381172
rect 262876 381108 262877 381172
rect 262811 381107 262877 381108
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 261234 298894 261854 334338
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 261234 262894 261854 298338
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 226894 261854 262338
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 190894 261854 226338
rect 262259 211852 262325 211853
rect 262259 211788 262260 211852
rect 262324 211788 262325 211852
rect 262259 211787 262325 211788
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 259683 186964 259749 186965
rect 259683 186900 259684 186964
rect 259748 186900 259749 186964
rect 259683 186899 259749 186900
rect 259686 158677 259746 186899
rect 259683 158676 259749 158677
rect 259683 158612 259684 158676
rect 259748 158612 259749 158676
rect 259683 158611 259749 158612
rect 261234 154894 261854 190338
rect 262075 175404 262141 175405
rect 262075 175340 262076 175404
rect 262140 175340 262141 175404
rect 262075 175339 262141 175340
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 262078 96661 262138 175339
rect 262262 161805 262322 211787
rect 262259 161804 262325 161805
rect 262259 161740 262260 161804
rect 262324 161740 262325 161804
rect 262259 161739 262325 161740
rect 262075 96660 262141 96661
rect 262075 96596 262076 96660
rect 262140 96596 262141 96660
rect 262075 96595 262141 96596
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 258395 3500 258461 3501
rect 258395 3436 258396 3500
rect 258460 3436 258461 3500
rect 258395 3435 258461 3436
rect 259499 3500 259565 3501
rect 259499 3436 259500 3500
rect 259564 3436 259565 3500
rect 259499 3435 259565 3436
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 -4186 261854 10338
rect 262814 3637 262874 381107
rect 264954 374614 265574 410058
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 273851 383756 273917 383757
rect 273851 383692 273852 383756
rect 273916 383692 273917 383756
rect 273851 383691 273917 383692
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 269619 368524 269685 368525
rect 269619 368460 269620 368524
rect 269684 368460 269685 368524
rect 269619 368459 269685 368460
rect 267779 364988 267845 364989
rect 267779 364924 267780 364988
rect 267844 364924 267845 364988
rect 267779 364923 267845 364924
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 263547 330444 263613 330445
rect 263547 330380 263548 330444
rect 263612 330380 263613 330444
rect 263547 330379 263613 330380
rect 262811 3636 262877 3637
rect 262811 3572 262812 3636
rect 262876 3572 262877 3636
rect 262811 3571 262877 3572
rect 263550 3501 263610 330379
rect 264954 302614 265574 338058
rect 266307 334660 266373 334661
rect 266307 334596 266308 334660
rect 266372 334596 266373 334660
rect 266307 334595 266373 334596
rect 265755 313988 265821 313989
rect 265755 313924 265756 313988
rect 265820 313924 265821 313988
rect 265755 313923 265821 313924
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 266614 265574 302058
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 230614 265574 266058
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 263731 176356 263797 176357
rect 263731 176292 263732 176356
rect 263796 176292 263797 176356
rect 263731 176291 263797 176292
rect 263734 157181 263794 176291
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 263731 157180 263797 157181
rect 263731 157116 263732 157180
rect 263796 157116 263797 157180
rect 263731 157115 263797 157116
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 263547 3500 263613 3501
rect 263547 3436 263548 3500
rect 263612 3436 263613 3500
rect 263547 3435 263613 3436
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 265758 3501 265818 313923
rect 266310 3501 266370 334595
rect 266491 178804 266557 178805
rect 266491 178740 266492 178804
rect 266556 178740 266557 178804
rect 266491 178739 266557 178740
rect 266494 141133 266554 178739
rect 266491 141132 266557 141133
rect 266491 141068 266492 141132
rect 266556 141068 266557 141132
rect 266491 141067 266557 141068
rect 267782 3637 267842 364923
rect 269622 14517 269682 368459
rect 271091 353564 271157 353565
rect 271091 353500 271092 353564
rect 271156 353500 271157 353564
rect 271091 353499 271157 353500
rect 271094 33829 271154 353499
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271091 33828 271157 33829
rect 271091 33764 271092 33828
rect 271156 33764 271157 33828
rect 271091 33763 271157 33764
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 269619 14516 269685 14517
rect 269619 14452 269620 14516
rect 269684 14452 269685 14516
rect 269619 14451 269685 14452
rect 267779 3636 267845 3637
rect 267779 3572 267780 3636
rect 267844 3572 267845 3636
rect 267779 3571 267845 3572
rect 265755 3500 265821 3501
rect 265755 3436 265756 3500
rect 265820 3436 265821 3500
rect 265755 3435 265821 3436
rect 266307 3500 266373 3501
rect 266307 3436 266308 3500
rect 266372 3436 266373 3500
rect 266307 3435 266373 3436
rect 271794 -1306 272414 20898
rect 273854 3365 273914 383691
rect 275514 349174 276134 384618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 276243 358052 276309 358053
rect 276243 357988 276244 358052
rect 276308 357988 276309 358052
rect 276243 357987 276309 357988
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 277174 276134 312618
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 205174 276134 240618
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 169174 276134 204618
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 133174 276134 168618
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 273851 3364 273917 3365
rect 273851 3300 273852 3364
rect 273916 3300 273917 3364
rect 273851 3299 273917 3300
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 -3226 276134 24618
rect 276246 3637 276306 357987
rect 279234 352894 279854 388338
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 280894 279854 316338
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279234 172894 279854 208338
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 279234 136894 279854 172338
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 100894 279854 136338
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 276243 3636 276309 3637
rect 276243 3572 276244 3636
rect 276308 3572 276309 3636
rect 276243 3571 276309 3572
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 356614 283574 392058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 286179 381036 286245 381037
rect 286179 380972 286180 381036
rect 286244 380972 286245 381036
rect 286179 380971 286245 380972
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 282954 284614 283574 320058
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 282954 248614 283574 284058
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 282954 176614 283574 212058
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 286182 3637 286242 380971
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 288387 325140 288453 325141
rect 288387 325076 288388 325140
rect 288452 325076 288453 325140
rect 288387 325075 288453 325076
rect 286179 3636 286245 3637
rect 286179 3572 286180 3636
rect 286244 3572 286245 3636
rect 286179 3571 286245 3572
rect 288390 3501 288450 325075
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 288387 3500 288453 3501
rect 288387 3436 288388 3500
rect 288452 3436 288453 3500
rect 288387 3435 288453 3436
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 298691 379540 298757 379541
rect 298691 379476 298692 379540
rect 298756 379476 298757 379540
rect 298691 379475 298757 379476
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 298694 3637 298754 379475
rect 300954 374614 301574 410058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 303659 380220 303725 380221
rect 303659 380156 303660 380220
rect 303724 380156 303725 380220
rect 303659 380155 303725 380156
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 301819 352612 301885 352613
rect 301819 352548 301820 352612
rect 301884 352548 301885 352612
rect 301819 352547 301885 352548
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 299979 113932 300045 113933
rect 299979 113868 299980 113932
rect 300044 113868 300045 113932
rect 299979 113867 300045 113868
rect 299982 53141 300042 113867
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 299979 53140 300045 53141
rect 299979 53076 299980 53140
rect 300044 53076 300045 53140
rect 299979 53075 300045 53076
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 298691 3636 298757 3637
rect 298691 3572 298692 3636
rect 298756 3572 298757 3636
rect 298691 3571 298757 3572
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 301822 3501 301882 352547
rect 302187 305692 302253 305693
rect 302187 305628 302188 305692
rect 302252 305628 302253 305692
rect 302187 305627 302253 305628
rect 302190 3501 302250 305627
rect 302739 139772 302805 139773
rect 302739 139708 302740 139772
rect 302804 139708 302805 139772
rect 302739 139707 302805 139708
rect 302742 36549 302802 139707
rect 302739 36548 302805 36549
rect 302739 36484 302740 36548
rect 302804 36484 302805 36548
rect 302739 36483 302805 36484
rect 303662 3501 303722 380155
rect 304947 377772 305013 377773
rect 304947 377708 304948 377772
rect 305012 377708 305013 377772
rect 304947 377707 305013 377708
rect 304211 131476 304277 131477
rect 304211 131412 304212 131476
rect 304276 131412 304277 131476
rect 304211 131411 304277 131412
rect 304214 64157 304274 131411
rect 304211 64156 304277 64157
rect 304211 64092 304212 64156
rect 304276 64092 304277 64156
rect 304211 64091 304277 64092
rect 304950 3501 305010 377707
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 178000 308414 200898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 178000 312134 204618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 178000 315854 208338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 321507 296852 321573 296853
rect 321507 296788 321508 296852
rect 321572 296788 321573 296852
rect 321507 296787 321573 296788
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 178000 319574 212058
rect 306971 175268 307037 175269
rect 306971 175204 306972 175268
rect 307036 175204 307037 175268
rect 306971 175203 307037 175204
rect 306974 141405 307034 175203
rect 314208 165454 314528 165486
rect 314208 165218 314250 165454
rect 314486 165218 314528 165454
rect 314208 165134 314528 165218
rect 314208 164898 314250 165134
rect 314486 164898 314528 165134
rect 314208 164866 314528 164898
rect 317472 165454 317792 165486
rect 317472 165218 317514 165454
rect 317750 165218 317792 165454
rect 317472 165134 317792 165218
rect 317472 164898 317514 165134
rect 317750 164898 317792 165134
rect 317472 164866 317792 164898
rect 312576 147454 312896 147486
rect 312576 147218 312618 147454
rect 312854 147218 312896 147454
rect 312576 147134 312896 147218
rect 312576 146898 312618 147134
rect 312854 146898 312896 147134
rect 312576 146866 312896 146898
rect 315840 147454 316160 147486
rect 315840 147218 315882 147454
rect 316118 147218 316160 147454
rect 315840 147134 316160 147218
rect 315840 146898 315882 147134
rect 316118 146898 316160 147134
rect 315840 146866 316160 146898
rect 319104 147454 319424 147486
rect 319104 147218 319146 147454
rect 319382 147218 319424 147454
rect 319104 147134 319424 147218
rect 319104 146898 319146 147134
rect 319382 146898 319424 147134
rect 319104 146866 319424 146898
rect 306971 141404 307037 141405
rect 306971 141340 306972 141404
rect 307036 141340 307037 141404
rect 306971 141339 307037 141340
rect 307523 141268 307589 141269
rect 307523 141204 307524 141268
rect 307588 141204 307589 141268
rect 307523 141203 307589 141204
rect 307526 131749 307586 141203
rect 321510 134469 321570 296787
rect 322979 293996 323045 293997
rect 322979 293932 322980 293996
rect 323044 293932 323045 293996
rect 322979 293931 323045 293932
rect 321507 134468 321573 134469
rect 321507 134404 321508 134468
rect 321572 134404 321573 134468
rect 321507 134403 321573 134404
rect 307523 131748 307589 131749
rect 307523 131684 307524 131748
rect 307588 131684 307589 131748
rect 307523 131683 307589 131684
rect 305499 130116 305565 130117
rect 305499 130052 305500 130116
rect 305564 130052 305565 130116
rect 305499 130051 305565 130052
rect 305502 62797 305562 130051
rect 314208 129454 314528 129486
rect 314208 129218 314250 129454
rect 314486 129218 314528 129454
rect 314208 129134 314528 129218
rect 314208 128898 314250 129134
rect 314486 128898 314528 129134
rect 314208 128866 314528 128898
rect 317472 129454 317792 129486
rect 317472 129218 317514 129454
rect 317750 129218 317792 129454
rect 317472 129134 317792 129218
rect 317472 128898 317514 129134
rect 317750 128898 317792 129134
rect 317472 128866 317792 128898
rect 306971 126444 307037 126445
rect 306971 126380 306972 126444
rect 307036 126380 307037 126444
rect 306971 126379 307037 126380
rect 305499 62796 305565 62797
rect 305499 62732 305500 62796
rect 305564 62732 305565 62796
rect 305499 62731 305565 62732
rect 306974 13021 307034 126379
rect 312576 111454 312896 111486
rect 312576 111218 312618 111454
rect 312854 111218 312896 111454
rect 312576 111134 312896 111218
rect 312576 110898 312618 111134
rect 312854 110898 312896 111134
rect 312576 110866 312896 110898
rect 315840 111454 316160 111486
rect 315840 111218 315882 111454
rect 316118 111218 316160 111454
rect 315840 111134 316160 111218
rect 315840 110898 315882 111134
rect 316118 110898 316160 111134
rect 315840 110866 316160 110898
rect 319104 111454 319424 111486
rect 319104 111218 319146 111454
rect 319382 111218 319424 111454
rect 319104 111134 319424 111218
rect 319104 110898 319146 111134
rect 319382 110898 319424 111134
rect 319104 110866 319424 110898
rect 322982 107133 323042 293931
rect 325794 291454 326414 326898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 331259 340100 331325 340101
rect 331259 340036 331260 340100
rect 331324 340036 331325 340100
rect 331259 340035 331325 340036
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 327027 291956 327093 291957
rect 327027 291892 327028 291956
rect 327092 291892 327093 291956
rect 327027 291891 327093 291892
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 327030 131749 327090 291891
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 328499 226948 328565 226949
rect 328499 226884 328500 226948
rect 328564 226884 328565 226948
rect 328499 226883 328565 226884
rect 327027 131748 327093 131749
rect 327027 131684 327028 131748
rect 327092 131684 327093 131748
rect 327027 131683 327093 131684
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 322979 107132 323045 107133
rect 322979 107068 322980 107132
rect 323044 107068 323045 107132
rect 322979 107067 323045 107068
rect 307155 97068 307221 97069
rect 307155 97004 307156 97068
rect 307220 97004 307221 97068
rect 307155 97003 307221 97004
rect 324451 97068 324517 97069
rect 324451 97004 324452 97068
rect 324516 97004 324517 97068
rect 324451 97003 324517 97004
rect 306971 13020 307037 13021
rect 306971 12956 306972 13020
rect 307036 12956 307037 13020
rect 306971 12955 307037 12956
rect 307158 4861 307218 97003
rect 307794 93454 308414 94000
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307155 4860 307221 4861
rect 307155 4796 307156 4860
rect 307220 4796 307221 4860
rect 307155 4795 307221 4796
rect 301819 3500 301885 3501
rect 301819 3436 301820 3500
rect 301884 3436 301885 3500
rect 301819 3435 301885 3436
rect 302187 3500 302253 3501
rect 302187 3436 302188 3500
rect 302252 3436 302253 3500
rect 302187 3435 302253 3436
rect 303659 3500 303725 3501
rect 303659 3436 303660 3500
rect 303724 3436 303725 3500
rect 303659 3435 303725 3436
rect 304947 3500 305013 3501
rect 304947 3436 304948 3500
rect 305012 3436 305013 3500
rect 304947 3435 305013 3436
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 61174 312134 94000
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 64894 315854 94000
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 68614 319574 94000
rect 324454 93669 324514 97003
rect 324451 93668 324517 93669
rect 324451 93604 324452 93668
rect 324516 93604 324517 93668
rect 324451 93603 324517 93604
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 75454 326414 110898
rect 328502 106317 328562 226883
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 328499 106316 328565 106317
rect 328499 106252 328500 106316
rect 328564 106252 328565 106316
rect 328499 106251 328565 106252
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 331262 3501 331322 340035
rect 333234 334894 333854 370338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 335859 366348 335925 366349
rect 335859 366284 335860 366348
rect 335924 366284 335925 366348
rect 335859 366283 335925 366284
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 334019 304196 334085 304197
rect 334019 304132 334020 304196
rect 334084 304132 334085 304196
rect 334019 304131 334085 304132
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 332547 253196 332613 253197
rect 332547 253132 332548 253196
rect 332612 253132 332613 253196
rect 332547 253131 332613 253132
rect 331443 180164 331509 180165
rect 331443 180100 331444 180164
rect 331508 180100 331509 180164
rect 331443 180099 331509 180100
rect 331446 111077 331506 180099
rect 331443 111076 331509 111077
rect 331443 111012 331444 111076
rect 331508 111012 331509 111076
rect 331443 111011 331509 111012
rect 332550 3501 332610 253131
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 331259 3500 331325 3501
rect 331259 3436 331260 3500
rect 331324 3436 331325 3500
rect 331259 3435 331325 3436
rect 332547 3500 332613 3501
rect 332547 3436 332548 3500
rect 332612 3436 332613 3500
rect 332547 3435 332613 3436
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 -4186 333854 10338
rect 334022 3637 334082 304131
rect 335123 177444 335189 177445
rect 335123 177380 335124 177444
rect 335188 177380 335189 177444
rect 335123 177379 335189 177380
rect 334203 177308 334269 177309
rect 334203 177244 334204 177308
rect 334268 177244 334269 177308
rect 334203 177243 334269 177244
rect 334019 3636 334085 3637
rect 334019 3572 334020 3636
rect 334084 3572 334085 3636
rect 334019 3571 334085 3572
rect 334206 3501 334266 177243
rect 335126 4045 335186 177379
rect 335123 4044 335189 4045
rect 335123 3980 335124 4044
rect 335188 3980 335189 4044
rect 335123 3979 335189 3980
rect 335862 3501 335922 366283
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 338251 331804 338317 331805
rect 338251 331740 338252 331804
rect 338316 331740 338317 331804
rect 338251 331739 338317 331740
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336779 206276 336845 206277
rect 336779 206212 336780 206276
rect 336844 206212 336845 206276
rect 336779 206211 336845 206212
rect 336782 115973 336842 206211
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 338254 180810 338314 331739
rect 339539 327724 339605 327725
rect 339539 327660 339540 327724
rect 339604 327660 339605 327724
rect 339539 327659 339605 327660
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336779 115972 336845 115973
rect 336779 115908 336780 115972
rect 336844 115908 336845 115972
rect 336779 115907 336845 115908
rect 336954 86614 337574 122058
rect 338070 180750 338314 180810
rect 338070 93870 338130 180750
rect 338251 180028 338317 180029
rect 338251 179964 338252 180028
rect 338316 179964 338317 180028
rect 338251 179963 338317 179964
rect 338254 101013 338314 179963
rect 338251 101012 338317 101013
rect 338251 100948 338252 101012
rect 338316 100948 338317 101012
rect 338251 100947 338317 100948
rect 338070 93810 338314 93870
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 334203 3500 334269 3501
rect 334203 3436 334204 3500
rect 334268 3436 334269 3500
rect 334203 3435 334269 3436
rect 335859 3500 335925 3501
rect 335859 3436 335860 3500
rect 335924 3436 335925 3500
rect 335859 3435 335925 3436
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 338254 3501 338314 93810
rect 339542 3501 339602 327659
rect 342299 325004 342365 325005
rect 342299 324940 342300 325004
rect 342364 324940 342365 325004
rect 342299 324939 342365 324940
rect 340827 319428 340893 319429
rect 340827 319364 340828 319428
rect 340892 319364 340893 319428
rect 340827 319363 340893 319364
rect 339723 192540 339789 192541
rect 339723 192476 339724 192540
rect 339788 192476 339789 192540
rect 339723 192475 339789 192476
rect 339726 124269 339786 192475
rect 339723 124268 339789 124269
rect 339723 124204 339724 124268
rect 339788 124204 339789 124268
rect 339723 124203 339789 124204
rect 340830 3501 340890 319363
rect 342302 3501 342362 324939
rect 343794 309454 344414 344898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 345059 309772 345125 309773
rect 345059 309708 345060 309772
rect 345124 309708 345125 309772
rect 345059 309707 345125 309708
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 338251 3500 338317 3501
rect 338251 3436 338252 3500
rect 338316 3436 338317 3500
rect 338251 3435 338317 3436
rect 339539 3500 339605 3501
rect 339539 3436 339540 3500
rect 339604 3436 339605 3500
rect 339539 3435 339605 3436
rect 340827 3500 340893 3501
rect 340827 3436 340828 3500
rect 340892 3436 340893 3500
rect 340827 3435 340893 3436
rect 342299 3500 342365 3501
rect 342299 3436 342300 3500
rect 342364 3436 342365 3500
rect 342299 3435 342365 3436
rect 343794 -1306 344414 20898
rect 345062 3501 345122 309707
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 345059 3500 345125 3501
rect 345059 3436 345060 3500
rect 345124 3436 345125 3500
rect 345059 3435 345125 3436
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 580211 282164 580277 282165
rect 580211 282100 580212 282164
rect 580276 282100 580277 282164
rect 580211 282099 580277 282100
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 580214 139365 580274 282099
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 580211 139364 580277 139365
rect 580211 139300 580212 139364
rect 580276 139300 580277 139364
rect 580211 139299 580277 139300
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 74250 363218 74486 363454
rect 74250 362898 74486 363134
rect 104970 363218 105206 363454
rect 104970 362898 105206 363134
rect 89610 345218 89846 345454
rect 89610 344898 89846 345134
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 89610 273218 89846 273454
rect 89610 272898 89846 273134
rect 74250 255218 74486 255454
rect 74250 254898 74486 255134
rect 104970 255218 105206 255454
rect 104970 254898 105206 255134
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 69128 165218 69364 165454
rect 69128 164898 69364 165134
rect 164192 165218 164428 165454
rect 164192 164898 164428 165134
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 69808 147218 70044 147454
rect 69808 146898 70044 147134
rect 163512 147218 163748 147454
rect 163512 146898 163748 147134
rect 69128 129218 69364 129454
rect 69128 128898 69364 129134
rect 164192 129218 164428 129454
rect 164192 128898 164428 129134
rect 69808 111218 70044 111454
rect 69808 110898 70044 111134
rect 163512 111218 163748 111454
rect 163512 110898 163748 111134
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 203546 276938 203782 277174
rect 203866 276938 204102 277174
rect 203546 276618 203782 276854
rect 203866 276618 204102 276854
rect 203546 240938 203782 241174
rect 203866 240938 204102 241174
rect 203546 240618 203782 240854
rect 203866 240618 204102 240854
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 207266 280658 207502 280894
rect 207586 280658 207822 280894
rect 207266 280338 207502 280574
rect 207586 280338 207822 280574
rect 207266 244658 207502 244894
rect 207586 244658 207822 244894
rect 207266 244338 207502 244574
rect 207586 244338 207822 244574
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 210986 284378 211222 284614
rect 211306 284378 211542 284614
rect 210986 284058 211222 284294
rect 211306 284058 211542 284294
rect 210986 248378 211222 248614
rect 211306 248378 211542 248614
rect 210986 248058 211222 248294
rect 211306 248058 211542 248294
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 239546 276938 239782 277174
rect 239866 276938 240102 277174
rect 239546 276618 239782 276854
rect 239866 276618 240102 276854
rect 239546 240938 239782 241174
rect 239866 240938 240102 241174
rect 239546 240618 239782 240854
rect 239866 240618 240102 240854
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 243266 280658 243502 280894
rect 243586 280658 243822 280894
rect 243266 280338 243502 280574
rect 243586 280338 243822 280574
rect 243266 244658 243502 244894
rect 243586 244658 243822 244894
rect 243266 244338 243502 244574
rect 243586 244338 243822 244574
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 246986 284378 247222 284614
rect 247306 284378 247542 284614
rect 246986 284058 247222 284294
rect 247306 284058 247542 284294
rect 246986 248378 247222 248614
rect 247306 248378 247542 248614
rect 246986 248058 247222 248294
rect 247306 248058 247542 248294
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 227916 165218 228152 165454
rect 227916 164898 228152 165134
rect 237847 165218 238083 165454
rect 237847 164898 238083 165134
rect 222952 147218 223188 147454
rect 222952 146898 223188 147134
rect 232882 147218 233118 147454
rect 232882 146898 233118 147134
rect 242813 147218 243049 147454
rect 242813 146898 243049 147134
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 227916 129218 228152 129454
rect 227916 128898 228152 129134
rect 237847 129218 238083 129454
rect 237847 128898 238083 129134
rect 222952 111218 223188 111454
rect 222952 110898 223188 111134
rect 232882 111218 233118 111454
rect 232882 110898 233118 111134
rect 242813 111218 243049 111454
rect 242813 110898 243049 111134
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 314250 165218 314486 165454
rect 314250 164898 314486 165134
rect 317514 165218 317750 165454
rect 317514 164898 317750 165134
rect 312618 147218 312854 147454
rect 312618 146898 312854 147134
rect 315882 147218 316118 147454
rect 315882 146898 316118 147134
rect 319146 147218 319382 147454
rect 319146 146898 319382 147134
rect 314250 129218 314486 129454
rect 314250 128898 314486 129134
rect 317514 129218 317750 129454
rect 317514 128898 317750 129134
rect 312618 111218 312854 111454
rect 312618 110898 312854 111134
rect 315882 111218 316118 111454
rect 315882 110898 316118 111134
rect 319146 111218 319382 111454
rect 319146 110898 319382 111134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 74250 363454
rect 74486 363218 104970 363454
rect 105206 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 74250 363134
rect 74486 362898 104970 363134
rect 105206 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 89610 345454
rect 89846 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 89610 345134
rect 89846 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 89610 273454
rect 89846 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 89610 273134
rect 89846 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 74250 255454
rect 74486 255218 104970 255454
rect 105206 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 74250 255134
rect 74486 254898 104970 255134
rect 105206 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 69128 165454
rect 69364 165218 164192 165454
rect 164428 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 227916 165454
rect 228152 165218 237847 165454
rect 238083 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 314250 165454
rect 314486 165218 317514 165454
rect 317750 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 69128 165134
rect 69364 164898 164192 165134
rect 164428 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 227916 165134
rect 228152 164898 237847 165134
rect 238083 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 314250 165134
rect 314486 164898 317514 165134
rect 317750 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 69808 147454
rect 70044 147218 163512 147454
rect 163748 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 222952 147454
rect 223188 147218 232882 147454
rect 233118 147218 242813 147454
rect 243049 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 312618 147454
rect 312854 147218 315882 147454
rect 316118 147218 319146 147454
rect 319382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 69808 147134
rect 70044 146898 163512 147134
rect 163748 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 222952 147134
rect 223188 146898 232882 147134
rect 233118 146898 242813 147134
rect 243049 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 312618 147134
rect 312854 146898 315882 147134
rect 316118 146898 319146 147134
rect 319382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 69128 129454
rect 69364 129218 164192 129454
rect 164428 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 227916 129454
rect 228152 129218 237847 129454
rect 238083 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 314250 129454
rect 314486 129218 317514 129454
rect 317750 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 69128 129134
rect 69364 128898 164192 129134
rect 164428 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 227916 129134
rect 228152 128898 237847 129134
rect 238083 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 314250 129134
rect 314486 128898 317514 129134
rect 317750 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 69808 111454
rect 70044 111218 163512 111454
rect 163748 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 222952 111454
rect 223188 111218 232882 111454
rect 233118 111218 242813 111454
rect 243049 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 312618 111454
rect 312854 111218 315882 111454
rect 316118 111218 319146 111454
rect 319382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 69808 111134
rect 70044 110898 163512 111134
rect 163748 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 222952 111134
rect 223188 110898 232882 111134
rect 233118 110898 242813 111134
rect 243049 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 312618 111134
rect 312854 110898 315882 111134
rect 316118 110898 319146 111134
rect 319382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_1kbyte_1rw1r_32x256_8  openram_1kB
timestamp 0
transform 1 0 68800 0 1 95100
box 0 0 95956 79500
use wb_bridge_2way  wb_bridge_2way
timestamp 0
transform 1 0 310000 0 1 96000
box 0 144 12000 80000
use wb_openram_wrapper  wb_openram_wrapper
timestamp 0
transform 1 0 217000 0 1 96000
box 0 144 32000 79688
use wrapped_cpr  wrapped_cpr_12
timestamp 0
transform 1 0 70000 0 1 340000
box -10 -52 40000 40000
use wrapped_function_generator  wrapped_function_generator_0
timestamp 0
transform 1 0 70000 0 1 240000
box 0 0 50000 52000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 94000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 176600 74414 238000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 176600 110414 238000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 294000 74414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 294000 110414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 382000 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 382000 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 176600 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 178000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 94000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 176600 78134 238000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 176600 114134 238000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 294000 78134 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 382000 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 294000 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 176600 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 178000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 94000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 176600 81854 238000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 176600 117854 238000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 294000 81854 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 382000 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 294000 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 176600 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 178000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 94000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 176600 85574 238000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 176600 121574 238000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 294000 85574 338000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 382000 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 294000 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 176600 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 178000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 94000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 94000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 176600 99854 238000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 294000 99854 338000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 382000 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 176600 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 178000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 178000 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 94000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 94000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 176600 103574 238000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 294000 103574 338000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 176600 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 382000 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 176600 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 178000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 178000 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 94000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 94000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 176600 92414 238000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 294000 92414 338000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 382000 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 176600 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 176600 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 178000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 178000 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 94000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 94000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 176600 96134 238000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 294000 96134 338000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 382000 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 176600 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 178000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 178000 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
