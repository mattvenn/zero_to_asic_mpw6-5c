magic
tech sky130A
magscale 1 2
timestamp 1650970008
<< metal1 >>
rect 201494 703060 201500 703112
rect 201552 703100 201558 703112
rect 202782 703100 202788 703112
rect 201552 703072 202788 703100
rect 201552 703060 201558 703072
rect 202782 703060 202788 703072
rect 202840 703060 202846 703112
rect 305638 703060 305644 703112
rect 305696 703100 305702 703112
rect 494790 703100 494796 703112
rect 305696 703072 494796 703100
rect 305696 703060 305702 703072
rect 494790 703060 494796 703072
rect 494848 703060 494854 703112
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 87598 702992 87604 703044
rect 87656 703032 87662 703044
rect 348786 703032 348792 703044
rect 87656 703004 348792 703032
rect 87656 702992 87662 703004
rect 348786 702992 348792 703004
rect 348844 702992 348850 703044
rect 107654 702924 107660 702976
rect 107712 702964 107718 702976
rect 413646 702964 413652 702976
rect 107712 702936 413652 702964
rect 107712 702924 107718 702936
rect 413646 702924 413652 702936
rect 413704 702924 413710 702976
rect 128998 702856 129004 702908
rect 129056 702896 129062 702908
rect 462314 702896 462320 702908
rect 129056 702868 462320 702896
rect 129056 702856 129062 702868
rect 462314 702856 462320 702868
rect 462372 702856 462378 702908
rect 53742 702788 53748 702840
rect 53800 702828 53806 702840
rect 397454 702828 397460 702840
rect 53800 702800 397460 702828
rect 53800 702788 53806 702800
rect 397454 702788 397460 702800
rect 397512 702788 397518 702840
rect 106274 702720 106280 702772
rect 106332 702760 106338 702772
rect 478506 702760 478512 702772
rect 106332 702732 478512 702760
rect 106332 702720 106338 702732
rect 478506 702720 478512 702732
rect 478564 702720 478570 702772
rect 57882 702652 57888 702704
rect 57940 702692 57946 702704
rect 429838 702692 429844 702704
rect 57940 702664 429844 702692
rect 57940 702652 57946 702664
rect 429838 702652 429844 702664
rect 429896 702652 429902 702704
rect 124858 702584 124864 702636
rect 124916 702624 124922 702636
rect 527174 702624 527180 702636
rect 124916 702596 527180 702624
rect 124916 702584 124922 702596
rect 527174 702584 527180 702596
rect 527232 702584 527238 702636
rect 133138 702516 133144 702568
rect 133196 702556 133202 702568
rect 559650 702556 559656 702568
rect 133196 702528 559656 702556
rect 133196 702516 133202 702528
rect 559650 702516 559656 702528
rect 559708 702516 559714 702568
rect 79318 702448 79324 702500
rect 79376 702488 79382 702500
rect 580902 702488 580908 702500
rect 79376 702460 580908 702488
rect 79376 702448 79382 702460
rect 580902 702448 580908 702460
rect 580960 702448 580966 702500
rect 55122 700340 55128 700392
rect 55180 700380 55186 700392
rect 105446 700380 105452 700392
rect 55180 700352 105452 700380
rect 55180 700340 55186 700352
rect 105446 700340 105452 700352
rect 105504 700340 105510 700392
rect 75178 700272 75184 700324
rect 75236 700312 75242 700324
rect 154114 700312 154120 700324
rect 75236 700284 154120 700312
rect 75236 700272 75242 700284
rect 154114 700272 154120 700284
rect 154172 700272 154178 700324
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 25498 699700 25504 699712
rect 24360 699672 25504 699700
rect 24360 699660 24366 699672
rect 25498 699660 25504 699672
rect 25556 699660 25562 699712
rect 214558 699660 214564 699712
rect 214616 699700 214622 699712
rect 218974 699700 218980 699712
rect 214616 699672 218980 699700
rect 214616 699660 214622 699672
rect 218974 699660 218980 699672
rect 219032 699660 219038 699712
rect 359458 699660 359464 699712
rect 359516 699700 359522 699712
rect 364978 699700 364984 699712
rect 359516 699672 364984 699700
rect 359516 699660 359522 699672
rect 364978 699660 364984 699672
rect 365036 699660 365042 699712
rect 151078 698912 151084 698964
rect 151136 698952 151142 698964
rect 235166 698952 235172 698964
rect 151136 698924 235172 698952
rect 151136 698912 151142 698924
rect 235166 698912 235172 698924
rect 235224 698912 235230 698964
rect 62022 697620 62028 697672
rect 62080 697660 62086 697672
rect 137830 697660 137836 697672
rect 62080 697632 137836 697660
rect 62080 697620 62086 697632
rect 137830 697620 137836 697632
rect 137888 697620 137894 697672
rect 266354 697620 266360 697672
rect 266412 697660 266418 697672
rect 267642 697660 267648 697672
rect 266412 697632 267648 697660
rect 266412 697620 266418 697632
rect 267642 697620 267648 697632
rect 267700 697620 267706 697672
rect 134518 697552 134524 697604
rect 134576 697592 134582 697604
rect 283834 697592 283840 697604
rect 134576 697564 283840 697592
rect 134576 697552 134582 697564
rect 283834 697552 283840 697564
rect 283892 697552 283898 697604
rect 126238 683136 126244 683188
rect 126296 683176 126302 683188
rect 580166 683176 580172 683188
rect 126296 683148 580172 683176
rect 126296 683136 126302 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 32398 670732 32404 670744
rect 3568 670704 32404 670732
rect 3568 670692 3574 670704
rect 32398 670692 32404 670704
rect 32456 670692 32462 670744
rect 148318 670692 148324 670744
rect 148376 670732 148382 670744
rect 580166 670732 580172 670744
rect 148376 670704 580172 670732
rect 148376 670692 148382 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3510 656888 3516 656940
rect 3568 656928 3574 656940
rect 15838 656928 15844 656940
rect 3568 656900 15844 656928
rect 3568 656888 3574 656900
rect 15838 656888 15844 656900
rect 15896 656888 15902 656940
rect 123478 643084 123484 643136
rect 123536 643124 123542 643136
rect 580166 643124 580172 643136
rect 123536 643096 580172 643124
rect 123536 643084 123542 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3510 632068 3516 632120
rect 3568 632108 3574 632120
rect 21358 632108 21364 632120
rect 3568 632080 21364 632108
rect 3568 632068 3574 632080
rect 21358 632068 21364 632080
rect 21416 632068 21422 632120
rect 3510 618264 3516 618316
rect 3568 618304 3574 618316
rect 17218 618304 17224 618316
rect 3568 618276 17224 618304
rect 3568 618264 3574 618276
rect 17218 618264 17224 618276
rect 17276 618264 17282 618316
rect 130378 616836 130384 616888
rect 130436 616876 130442 616888
rect 580166 616876 580172 616888
rect 130436 616848 580172 616876
rect 130436 616836 130442 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3510 605820 3516 605872
rect 3568 605860 3574 605872
rect 14458 605860 14464 605872
rect 3568 605832 14464 605860
rect 3568 605820 3574 605832
rect 14458 605820 14464 605832
rect 14516 605820 14522 605872
rect 52362 590656 52368 590708
rect 52420 590696 52426 590708
rect 579798 590696 579804 590708
rect 52420 590668 579804 590696
rect 52420 590656 52426 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 116578 579680 116584 579692
rect 3384 579652 116584 579680
rect 3384 579640 3390 579652
rect 116578 579640 116584 579652
rect 116636 579640 116642 579692
rect 142798 576852 142804 576904
rect 142856 576892 142862 576904
rect 580166 576892 580172 576904
rect 142856 576864 580172 576892
rect 142856 576852 142862 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3234 565836 3240 565888
rect 3292 565876 3298 565888
rect 29638 565876 29644 565888
rect 3292 565848 29644 565876
rect 3292 565836 3298 565848
rect 29638 565836 29644 565848
rect 29696 565836 29702 565888
rect 97258 563048 97264 563100
rect 97316 563088 97322 563100
rect 579798 563088 579804 563100
rect 97316 563060 579804 563088
rect 97316 563048 97322 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 18598 553432 18604 553444
rect 3384 553404 18604 553432
rect 3384 553392 3390 553404
rect 18598 553392 18604 553404
rect 18656 553392 18662 553444
rect 123570 536800 123576 536852
rect 123628 536840 123634 536852
rect 580166 536840 580172 536852
rect 123628 536812 580172 536840
rect 123628 536800 123634 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 2958 527144 2964 527196
rect 3016 527184 3022 527196
rect 39298 527184 39304 527196
rect 3016 527156 39304 527184
rect 3016 527144 3022 527156
rect 39298 527144 39304 527156
rect 39356 527144 39362 527196
rect 141418 524424 141424 524476
rect 141476 524464 141482 524476
rect 580166 524464 580172 524476
rect 141476 524436 580172 524464
rect 141476 524424 141482 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 66162 510620 66168 510672
rect 66220 510660 66226 510672
rect 580166 510660 580172 510672
rect 66220 510632 580172 510660
rect 66220 510620 66226 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3326 500964 3332 501016
rect 3384 501004 3390 501016
rect 120074 501004 120080 501016
rect 3384 500976 120080 501004
rect 3384 500964 3390 500976
rect 120074 500964 120080 500976
rect 120132 500964 120138 501016
rect 126330 484372 126336 484424
rect 126388 484412 126394 484424
rect 580166 484412 580172 484424
rect 126388 484384 580172 484412
rect 126388 484372 126394 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 3050 474716 3056 474768
rect 3108 474756 3114 474768
rect 111058 474756 111064 474768
rect 3108 474728 111064 474756
rect 3108 474716 3114 474728
rect 111058 474716 111064 474728
rect 111116 474716 111122 474768
rect 124950 470568 124956 470620
rect 125008 470608 125014 470620
rect 579982 470608 579988 470620
rect 125008 470580 579988 470608
rect 125008 470568 125014 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3326 462340 3332 462392
rect 3384 462380 3390 462392
rect 47578 462380 47584 462392
rect 3384 462352 47584 462380
rect 3384 462340 3390 462352
rect 47578 462340 47584 462352
rect 47636 462340 47642 462392
rect 3326 448536 3332 448588
rect 3384 448576 3390 448588
rect 22738 448576 22744 448588
rect 3384 448548 22744 448576
rect 3384 448536 3390 448548
rect 22738 448536 22744 448548
rect 22796 448536 22802 448588
rect 129090 430584 129096 430636
rect 129148 430624 129154 430636
rect 580166 430624 580172 430636
rect 129148 430596 580172 430624
rect 129148 430584 129154 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 2774 423512 2780 423564
rect 2832 423552 2838 423564
rect 4798 423552 4804 423564
rect 2832 423524 4804 423552
rect 2832 423512 2838 423524
rect 4798 423512 4804 423524
rect 4856 423512 4862 423564
rect 93118 418140 93124 418192
rect 93176 418180 93182 418192
rect 580166 418180 580172 418192
rect 93176 418152 580172 418180
rect 93176 418140 93182 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 3326 409844 3332 409896
rect 3384 409884 3390 409896
rect 33778 409884 33784 409896
rect 3384 409856 33784 409884
rect 3384 409844 3390 409856
rect 33778 409844 33784 409856
rect 33836 409844 33842 409896
rect 67542 404336 67548 404388
rect 67600 404376 67606 404388
rect 580166 404376 580172 404388
rect 67600 404348 580172 404376
rect 67600 404336 67606 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3326 397468 3332 397520
rect 3384 397508 3390 397520
rect 35158 397508 35164 397520
rect 3384 397480 35164 397508
rect 3384 397468 3390 397480
rect 35158 397468 35164 397480
rect 35216 397468 35222 397520
rect 127618 378156 127624 378208
rect 127676 378196 127682 378208
rect 580166 378196 580172 378208
rect 127676 378168 580172 378196
rect 127676 378156 127682 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 3326 371220 3332 371272
rect 3384 371260 3390 371272
rect 43438 371260 43444 371272
rect 3384 371232 43444 371260
rect 3384 371220 3390 371232
rect 43438 371220 43444 371232
rect 43496 371220 43502 371272
rect 3326 357416 3332 357468
rect 3384 357456 3390 357468
rect 54478 357456 54484 357468
rect 3384 357428 54484 357456
rect 3384 357416 3390 357428
rect 54478 357416 54484 357428
rect 54536 357416 54542 357468
rect 76558 351908 76564 351960
rect 76616 351948 76622 351960
rect 580166 351948 580172 351960
rect 76616 351920 580172 351948
rect 76616 351908 76622 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 101398 345080 101404 345092
rect 3384 345052 101404 345080
rect 3384 345040 3390 345052
rect 101398 345040 101404 345052
rect 101456 345040 101462 345092
rect 88334 327700 88340 327752
rect 88392 327740 88398 327752
rect 103790 327740 103796 327752
rect 88392 327712 103796 327740
rect 88392 327700 88398 327712
rect 103790 327700 103796 327712
rect 103848 327700 103854 327752
rect 3418 324912 3424 324964
rect 3476 324952 3482 324964
rect 120258 324952 120264 324964
rect 3476 324924 120264 324952
rect 3476 324912 3482 324924
rect 120258 324912 120264 324924
rect 120316 324912 120322 324964
rect 91094 319404 91100 319456
rect 91152 319444 91158 319456
rect 148318 319444 148324 319456
rect 91152 319416 148324 319444
rect 91152 319404 91158 319416
rect 148318 319404 148324 319416
rect 148376 319404 148382 319456
rect 3326 318792 3332 318844
rect 3384 318832 3390 318844
rect 11698 318832 11704 318844
rect 3384 318804 11704 318832
rect 3384 318792 3390 318804
rect 11698 318792 11704 318804
rect 11756 318792 11762 318844
rect 116578 318724 116584 318776
rect 116636 318764 116642 318776
rect 121454 318764 121460 318776
rect 116636 318736 121460 318764
rect 116636 318724 116642 318736
rect 121454 318724 121460 318736
rect 121512 318724 121518 318776
rect 11698 318044 11704 318096
rect 11756 318084 11762 318096
rect 115934 318084 115940 318096
rect 11756 318056 115940 318084
rect 11756 318044 11762 318056
rect 115934 318044 115940 318056
rect 115992 318044 115998 318096
rect 93946 317500 93952 317552
rect 94004 317540 94010 317552
rect 97258 317540 97264 317552
rect 94004 317512 97264 317540
rect 94004 317500 94010 317512
rect 97258 317500 97264 317512
rect 97316 317500 97322 317552
rect 3510 315256 3516 315308
rect 3568 315296 3574 315308
rect 120166 315296 120172 315308
rect 3568 315268 120172 315296
rect 3568 315256 3574 315268
rect 120166 315256 120172 315268
rect 120224 315256 120230 315308
rect 77294 313896 77300 313948
rect 77352 313936 77358 313948
rect 93118 313936 93124 313948
rect 77352 313908 93124 313936
rect 77352 313896 77358 313908
rect 93118 313896 93124 313908
rect 93176 313896 93182 313948
rect 54478 312536 54484 312588
rect 54536 312576 54542 312588
rect 97994 312576 98000 312588
rect 54536 312548 98000 312576
rect 54536 312536 54542 312548
rect 97994 312536 98000 312548
rect 98052 312536 98058 312588
rect 125042 312536 125048 312588
rect 125100 312576 125106 312588
rect 580258 312576 580264 312588
rect 125100 312548 580264 312576
rect 125100 312536 125106 312548
rect 580258 312536 580264 312548
rect 580316 312536 580322 312588
rect 14458 311108 14464 311160
rect 14516 311148 14522 311160
rect 94130 311148 94136 311160
rect 14516 311120 94136 311148
rect 14516 311108 14522 311120
rect 94130 311108 94136 311120
rect 94188 311108 94194 311160
rect 101398 311108 101404 311160
rect 101456 311148 101462 311160
rect 118694 311148 118700 311160
rect 101456 311120 118700 311148
rect 101456 311108 101462 311120
rect 118694 311108 118700 311120
rect 118752 311108 118758 311160
rect 15838 309748 15844 309800
rect 15896 309788 15902 309800
rect 121546 309788 121552 309800
rect 15896 309760 121552 309788
rect 15896 309748 15902 309760
rect 121546 309748 121552 309760
rect 121604 309748 121610 309800
rect 123662 309748 123668 309800
rect 123720 309788 123726 309800
rect 580166 309788 580172 309800
rect 123720 309760 580172 309788
rect 123720 309748 123726 309760
rect 580166 309748 580172 309760
rect 580224 309748 580230 309800
rect 71774 308388 71780 308440
rect 71832 308428 71838 308440
rect 114554 308428 114560 308440
rect 71832 308400 114560 308428
rect 71832 308388 71838 308400
rect 114554 308388 114560 308400
rect 114612 308388 114618 308440
rect 122098 308388 122104 308440
rect 122156 308428 122162 308440
rect 201494 308428 201500 308440
rect 122156 308400 201500 308428
rect 122156 308388 122162 308400
rect 201494 308388 201500 308400
rect 201552 308388 201558 308440
rect 63402 307776 63408 307828
rect 63460 307816 63466 307828
rect 286318 307816 286324 307828
rect 63460 307788 286324 307816
rect 63460 307776 63466 307788
rect 286318 307776 286324 307788
rect 286376 307776 286382 307828
rect 89714 306348 89720 306400
rect 89772 306388 89778 306400
rect 302878 306388 302884 306400
rect 89772 306360 302884 306388
rect 89772 306348 89778 306360
rect 302878 306348 302884 306360
rect 302936 306348 302942 306400
rect 69014 305600 69020 305652
rect 69072 305640 69078 305652
rect 169754 305640 169760 305652
rect 69072 305612 169760 305640
rect 69072 305600 69078 305612
rect 169754 305600 169760 305612
rect 169812 305600 169818 305652
rect 92658 305056 92664 305108
rect 92716 305096 92722 305108
rect 233878 305096 233884 305108
rect 92716 305068 233884 305096
rect 92716 305056 92722 305068
rect 233878 305056 233884 305068
rect 233936 305056 233942 305108
rect 3234 304988 3240 305040
rect 3292 305028 3298 305040
rect 70394 305028 70400 305040
rect 3292 305000 70400 305028
rect 3292 304988 3298 305000
rect 70394 304988 70400 305000
rect 70452 304988 70458 305040
rect 75914 304988 75920 305040
rect 75972 305028 75978 305040
rect 287698 305028 287704 305040
rect 75972 305000 287704 305028
rect 75972 304988 75978 305000
rect 287698 304988 287704 305000
rect 287756 304988 287762 305040
rect 25498 304240 25504 304292
rect 25556 304280 25562 304292
rect 84470 304280 84476 304292
rect 25556 304252 84476 304280
rect 25556 304240 25562 304252
rect 84470 304240 84476 304252
rect 84528 304240 84534 304292
rect 85574 303764 85580 303816
rect 85632 303804 85638 303816
rect 170398 303804 170404 303816
rect 85632 303776 170404 303804
rect 85632 303764 85638 303776
rect 170398 303764 170404 303776
rect 170456 303764 170462 303816
rect 81894 303696 81900 303748
rect 81952 303736 81958 303748
rect 244918 303736 244924 303748
rect 81952 303708 244924 303736
rect 81952 303696 81958 303708
rect 244918 303696 244924 303708
rect 244976 303696 244982 303748
rect 74534 303628 74540 303680
rect 74592 303668 74598 303680
rect 267734 303668 267740 303680
rect 74592 303640 267740 303668
rect 74592 303628 74598 303640
rect 267734 303628 267740 303640
rect 267792 303628 267798 303680
rect 90358 302404 90364 302456
rect 90416 302444 90422 302456
rect 213178 302444 213184 302456
rect 90416 302416 213184 302444
rect 90416 302404 90422 302416
rect 213178 302404 213184 302416
rect 213236 302404 213242 302456
rect 69658 302336 69664 302388
rect 69716 302376 69722 302388
rect 224218 302376 224224 302388
rect 69716 302348 224224 302376
rect 69716 302336 69722 302348
rect 224218 302336 224224 302348
rect 224276 302336 224282 302388
rect 100846 302268 100852 302320
rect 100904 302308 100910 302320
rect 281534 302308 281540 302320
rect 100904 302280 281540 302308
rect 100904 302268 100910 302280
rect 281534 302268 281540 302280
rect 281592 302268 281598 302320
rect 71774 302200 71780 302252
rect 71832 302240 71838 302252
rect 334618 302240 334624 302252
rect 71832 302212 334624 302240
rect 71832 302200 71838 302212
rect 334618 302200 334624 302212
rect 334676 302200 334682 302252
rect 22738 301452 22744 301504
rect 22796 301492 22802 301504
rect 22796 301464 64874 301492
rect 22796 301452 22802 301464
rect 64846 301356 64874 301464
rect 70394 301452 70400 301504
rect 70452 301492 70458 301504
rect 121638 301492 121644 301504
rect 70452 301464 121644 301492
rect 70452 301452 70458 301464
rect 121638 301452 121644 301464
rect 121696 301452 121702 301504
rect 70394 301356 70400 301368
rect 64846 301328 70400 301356
rect 70394 301316 70400 301328
rect 70452 301316 70458 301368
rect 85666 300908 85672 300960
rect 85724 300948 85730 300960
rect 220078 300948 220084 300960
rect 85724 300920 220084 300948
rect 85724 300908 85730 300920
rect 220078 300908 220084 300920
rect 220136 300908 220142 300960
rect 102134 300840 102140 300892
rect 102192 300880 102198 300892
rect 280154 300880 280160 300892
rect 102192 300852 280160 300880
rect 102192 300840 102198 300852
rect 280154 300840 280160 300852
rect 280212 300840 280218 300892
rect 102318 299684 102324 299736
rect 102376 299724 102382 299736
rect 206278 299724 206284 299736
rect 102376 299696 206284 299724
rect 102376 299684 102382 299696
rect 206278 299684 206284 299696
rect 206336 299684 206342 299736
rect 84286 299616 84292 299668
rect 84344 299656 84350 299668
rect 202138 299656 202144 299668
rect 84344 299628 202144 299656
rect 84344 299616 84350 299628
rect 202138 299616 202144 299628
rect 202196 299616 202202 299668
rect 70486 299548 70492 299600
rect 70544 299588 70550 299600
rect 325786 299588 325792 299600
rect 70544 299560 325792 299588
rect 70544 299548 70550 299560
rect 325786 299548 325792 299560
rect 325844 299548 325850 299600
rect 80054 299480 80060 299532
rect 80112 299520 80118 299532
rect 583018 299520 583024 299532
rect 80112 299492 583024 299520
rect 80112 299480 80118 299492
rect 583018 299480 583024 299492
rect 583076 299480 583082 299532
rect 4798 298732 4804 298784
rect 4856 298772 4862 298784
rect 72602 298772 72608 298784
rect 4856 298744 72608 298772
rect 4856 298732 4862 298744
rect 72602 298732 72608 298744
rect 72660 298732 72666 298784
rect 89346 298460 89352 298512
rect 89404 298500 89410 298512
rect 148318 298500 148324 298512
rect 89404 298472 148324 298500
rect 89404 298460 89410 298472
rect 148318 298460 148324 298472
rect 148376 298460 148382 298512
rect 110598 298392 110604 298444
rect 110656 298432 110662 298444
rect 186958 298432 186964 298444
rect 110656 298404 186964 298432
rect 110656 298392 110662 298404
rect 186958 298392 186964 298404
rect 187016 298392 187022 298444
rect 79686 298324 79692 298376
rect 79744 298364 79750 298376
rect 197998 298364 198004 298376
rect 79744 298336 198004 298364
rect 79744 298324 79750 298336
rect 197998 298324 198004 298336
rect 198056 298324 198062 298376
rect 83550 298256 83556 298308
rect 83608 298296 83614 298308
rect 226978 298296 226984 298308
rect 83608 298268 226984 298296
rect 83608 298256 83614 298268
rect 226978 298256 226984 298268
rect 227036 298256 227042 298308
rect 111242 298188 111248 298240
rect 111300 298228 111306 298240
rect 345106 298228 345112 298240
rect 111300 298200 345112 298228
rect 111300 298188 111306 298200
rect 345106 298188 345112 298200
rect 345164 298188 345170 298240
rect 73890 298120 73896 298172
rect 73948 298160 73954 298172
rect 76558 298160 76564 298172
rect 73948 298132 76564 298160
rect 73948 298120 73954 298132
rect 76558 298120 76564 298132
rect 76616 298120 76622 298172
rect 88702 298120 88708 298172
rect 88760 298160 88766 298172
rect 335354 298160 335360 298172
rect 88760 298132 335360 298160
rect 88760 298120 88766 298132
rect 335354 298120 335360 298132
rect 335412 298120 335418 298172
rect 112530 297032 112536 297084
rect 112588 297072 112594 297084
rect 169018 297072 169024 297084
rect 112588 297044 169024 297072
rect 112588 297032 112594 297044
rect 169018 297032 169024 297044
rect 169076 297032 169082 297084
rect 82906 296964 82912 297016
rect 82964 297004 82970 297016
rect 215938 297004 215944 297016
rect 82964 296976 215944 297004
rect 82964 296964 82970 296976
rect 215938 296964 215944 296976
rect 215996 296964 216002 297016
rect 117682 296896 117688 296948
rect 117740 296936 117746 296948
rect 308398 296936 308404 296948
rect 117740 296908 308404 296936
rect 117740 296896 117746 296908
rect 308398 296896 308404 296908
rect 308456 296896 308462 296948
rect 113818 296828 113824 296880
rect 113876 296868 113882 296880
rect 346394 296868 346400 296880
rect 113876 296840 346400 296868
rect 113876 296828 113882 296840
rect 346394 296828 346400 296840
rect 346452 296828 346458 296880
rect 97718 296760 97724 296812
rect 97776 296800 97782 296812
rect 338114 296800 338120 296812
rect 97776 296772 338120 296800
rect 97776 296760 97782 296772
rect 338114 296760 338120 296772
rect 338172 296760 338178 296812
rect 77110 296692 77116 296744
rect 77168 296732 77174 296744
rect 342898 296732 342904 296744
rect 77168 296704 342904 296732
rect 77168 296692 77174 296704
rect 342898 296692 342904 296704
rect 342956 296692 342962 296744
rect 99650 295672 99656 295724
rect 99708 295712 99714 295724
rect 146938 295712 146944 295724
rect 99708 295684 146944 295712
rect 99708 295672 99714 295684
rect 146938 295672 146944 295684
rect 146996 295672 147002 295724
rect 11698 295604 11704 295656
rect 11756 295644 11762 295656
rect 118326 295644 118332 295656
rect 11756 295616 118332 295644
rect 11756 295604 11762 295616
rect 118326 295604 118332 295616
rect 118384 295604 118390 295656
rect 88058 295536 88064 295588
rect 88116 295576 88122 295588
rect 204898 295576 204904 295588
rect 88116 295548 204904 295576
rect 88116 295536 88122 295548
rect 204898 295536 204904 295548
rect 204956 295536 204962 295588
rect 68738 295468 68744 295520
rect 68796 295508 68802 295520
rect 252554 295508 252560 295520
rect 68796 295480 252560 295508
rect 68796 295468 68802 295480
rect 252554 295468 252560 295480
rect 252612 295468 252618 295520
rect 75178 295400 75184 295452
rect 75236 295440 75242 295452
rect 277394 295440 277400 295452
rect 75236 295412 277400 295440
rect 75236 295400 75242 295412
rect 277394 295400 277400 295412
rect 277452 295400 277458 295452
rect 99006 295332 99012 295384
rect 99064 295372 99070 295384
rect 336734 295372 336740 295384
rect 99064 295344 336740 295372
rect 99064 295332 99070 295344
rect 336734 295332 336740 295344
rect 336792 295332 336798 295384
rect 85482 295060 85488 295112
rect 85540 295100 85546 295112
rect 87598 295100 87604 295112
rect 85540 295072 87604 295100
rect 85540 295060 85546 295072
rect 87598 295060 87604 295072
rect 87656 295060 87662 295112
rect 73246 294584 73252 294636
rect 73304 294624 73310 294636
rect 111794 294624 111800 294636
rect 73304 294596 111800 294624
rect 73304 294584 73310 294596
rect 111794 294584 111800 294596
rect 111852 294584 111858 294636
rect 70394 294312 70400 294364
rect 70452 294352 70458 294364
rect 71038 294352 71044 294364
rect 70452 294324 71044 294352
rect 70452 294312 70458 294324
rect 71038 294312 71044 294324
rect 71096 294312 71102 294364
rect 77754 294312 77760 294364
rect 77812 294352 77818 294364
rect 79318 294352 79324 294364
rect 77812 294324 79324 294352
rect 77812 294312 77818 294324
rect 79318 294312 79324 294324
rect 79376 294312 79382 294364
rect 85574 294312 85580 294364
rect 85632 294352 85638 294364
rect 86494 294352 86500 294364
rect 85632 294324 86500 294352
rect 85632 294312 85638 294324
rect 86494 294312 86500 294324
rect 86552 294312 86558 294364
rect 93946 294312 93952 294364
rect 94004 294352 94010 294364
rect 94774 294352 94780 294364
rect 94004 294324 94780 294352
rect 94004 294312 94010 294324
rect 94774 294312 94780 294324
rect 94832 294312 94838 294364
rect 106734 294312 106740 294364
rect 106792 294352 106798 294364
rect 119706 294352 119712 294364
rect 106792 294324 119712 294352
rect 106792 294312 106798 294324
rect 119706 294312 119712 294324
rect 119764 294312 119770 294364
rect 67450 294244 67456 294296
rect 67508 294284 67514 294296
rect 92566 294284 92572 294296
rect 67508 294256 92572 294284
rect 67508 294244 67514 294256
rect 92566 294244 92572 294256
rect 92624 294244 92630 294296
rect 111886 294244 111892 294296
rect 111944 294284 111950 294296
rect 152458 294284 152464 294296
rect 111944 294256 152464 294284
rect 111944 294244 111950 294256
rect 152458 294244 152464 294256
rect 152516 294244 152522 294296
rect 87414 294176 87420 294228
rect 87472 294216 87478 294228
rect 137278 294216 137284 294228
rect 87472 294188 137284 294216
rect 87472 294176 87478 294188
rect 137278 294176 137284 294188
rect 137336 294176 137342 294228
rect 91922 294108 91928 294160
rect 91980 294148 91986 294160
rect 255406 294148 255412 294160
rect 91980 294120 255412 294148
rect 91980 294108 91986 294120
rect 255406 294108 255412 294120
rect 255464 294108 255470 294160
rect 3418 294040 3424 294092
rect 3476 294080 3482 294092
rect 97074 294080 97080 294092
rect 3476 294052 97080 294080
rect 3476 294040 3482 294052
rect 97074 294040 97080 294052
rect 97132 294040 97138 294092
rect 114462 294040 114468 294092
rect 114520 294080 114526 294092
rect 307018 294080 307024 294092
rect 114520 294052 307024 294080
rect 114520 294040 114526 294052
rect 307018 294040 307024 294052
rect 307076 294040 307082 294092
rect 50338 293972 50344 294024
rect 50396 294012 50402 294024
rect 79042 294012 79048 294024
rect 50396 293984 79048 294012
rect 50396 293972 50402 293984
rect 79042 293972 79048 293984
rect 79100 293972 79106 294024
rect 81618 293972 81624 294024
rect 81676 294012 81682 294024
rect 342254 294012 342260 294024
rect 81676 293984 342260 294012
rect 81676 293972 81682 293984
rect 342254 293972 342260 293984
rect 342312 293972 342318 294024
rect 111058 293224 111064 293276
rect 111116 293264 111122 293276
rect 125594 293264 125600 293276
rect 111116 293236 125600 293264
rect 111116 293224 111122 293236
rect 125594 293224 125600 293236
rect 125652 293224 125658 293276
rect 2774 292816 2780 292868
rect 2832 292856 2838 292868
rect 4798 292856 4804 292868
rect 2832 292828 4804 292856
rect 2832 292816 2838 292828
rect 4798 292816 4804 292828
rect 4856 292816 4862 292868
rect 8202 292816 8208 292868
rect 8260 292856 8266 292868
rect 96430 292856 96436 292868
rect 8260 292828 96436 292856
rect 8260 292816 8266 292828
rect 96430 292816 96436 292828
rect 96488 292816 96494 292868
rect 109310 292816 109316 292868
rect 109368 292856 109374 292868
rect 162118 292856 162124 292868
rect 109368 292828 162124 292856
rect 109368 292816 109374 292828
rect 162118 292816 162124 292828
rect 162176 292816 162182 292868
rect 53098 292748 53104 292800
rect 53156 292788 53162 292800
rect 101582 292788 101588 292800
rect 53156 292760 101588 292788
rect 53156 292748 53162 292760
rect 101582 292748 101588 292760
rect 101640 292748 101646 292800
rect 103514 292748 103520 292800
rect 103572 292788 103578 292800
rect 160738 292788 160744 292800
rect 103572 292760 160744 292788
rect 103572 292748 103578 292760
rect 160738 292748 160744 292760
rect 160796 292748 160802 292800
rect 93854 292680 93860 292732
rect 93912 292720 93918 292732
rect 178678 292720 178684 292732
rect 93912 292692 178684 292720
rect 93912 292680 93918 292692
rect 178678 292680 178684 292692
rect 178736 292680 178742 292732
rect 80974 292612 80980 292664
rect 81032 292652 81038 292664
rect 270494 292652 270500 292664
rect 81032 292624 270500 292652
rect 81032 292612 81038 292624
rect 270494 292612 270500 292624
rect 270552 292612 270558 292664
rect 68922 292544 68928 292596
rect 68980 292584 68986 292596
rect 267826 292584 267832 292596
rect 68980 292556 267832 292584
rect 68980 292544 68986 292556
rect 267826 292544 267832 292556
rect 267884 292544 267890 292596
rect 119062 291932 119068 291984
rect 119120 291972 119126 291984
rect 119798 291972 119804 291984
rect 119120 291944 119804 291972
rect 119120 291932 119126 291944
rect 119798 291932 119804 291944
rect 119856 291932 119862 291984
rect 115842 291864 115848 291916
rect 115900 291864 115906 291916
rect 117222 291864 117228 291916
rect 117280 291904 117286 291916
rect 117280 291876 122834 291904
rect 117280 291864 117286 291876
rect 3510 291796 3516 291848
rect 3568 291836 3574 291848
rect 67450 291836 67456 291848
rect 3568 291808 67456 291836
rect 3568 291796 3574 291808
rect 67450 291796 67456 291808
rect 67508 291796 67514 291848
rect 115860 291292 115888 291864
rect 122806 291360 122834 291876
rect 155218 291360 155224 291372
rect 122806 291332 155224 291360
rect 155218 291320 155224 291332
rect 155276 291320 155282 291372
rect 340874 291292 340880 291304
rect 115860 291264 340880 291292
rect 340874 291252 340880 291264
rect 340932 291252 340938 291304
rect 69750 291184 69756 291236
rect 69808 291224 69814 291236
rect 582742 291224 582748 291236
rect 69808 291196 582748 291224
rect 69808 291184 69814 291196
rect 582742 291184 582748 291196
rect 582800 291184 582806 291236
rect 121546 289892 121552 289944
rect 121604 289932 121610 289944
rect 255314 289932 255320 289944
rect 121604 289904 255320 289932
rect 121604 289892 121610 289904
rect 255314 289892 255320 289904
rect 255372 289892 255378 289944
rect 25498 289824 25504 289876
rect 25556 289864 25562 289876
rect 67634 289864 67640 289876
rect 25556 289836 67640 289864
rect 25556 289824 25562 289836
rect 67634 289824 67640 289836
rect 67692 289824 67698 289876
rect 121730 289824 121736 289876
rect 121788 289864 121794 289876
rect 269114 289864 269120 289876
rect 121788 289836 269120 289864
rect 121788 289824 121794 289836
rect 269114 289824 269120 289836
rect 269172 289824 269178 289876
rect 121546 289756 121552 289808
rect 121604 289796 121610 289808
rect 127618 289796 127624 289808
rect 121604 289768 127624 289796
rect 121604 289756 121610 289768
rect 127618 289756 127624 289768
rect 127676 289756 127682 289808
rect 121546 287036 121552 287088
rect 121604 287076 121610 287088
rect 351914 287076 351920 287088
rect 121604 287048 351920 287076
rect 121604 287036 121610 287048
rect 351914 287036 351920 287048
rect 351972 287036 351978 287088
rect 32398 286968 32404 287020
rect 32456 287008 32462 287020
rect 67634 287008 67640 287020
rect 32456 286980 67640 287008
rect 32456 286968 32462 286980
rect 67634 286968 67640 286980
rect 67692 286968 67698 287020
rect 122006 286288 122012 286340
rect 122064 286328 122070 286340
rect 329834 286328 329840 286340
rect 122064 286300 329840 286328
rect 122064 286288 122070 286300
rect 329834 286288 329840 286300
rect 329892 286288 329898 286340
rect 59078 285676 59084 285728
rect 59136 285716 59142 285728
rect 67726 285716 67732 285728
rect 59136 285688 67732 285716
rect 59136 285676 59142 285688
rect 67726 285676 67732 285688
rect 67784 285676 67790 285728
rect 63402 285608 63408 285660
rect 63460 285648 63466 285660
rect 67634 285648 67640 285660
rect 63460 285620 67640 285648
rect 63460 285608 63466 285620
rect 67634 285608 67640 285620
rect 67692 285608 67698 285660
rect 121638 285540 121644 285592
rect 121696 285580 121702 285592
rect 124950 285580 124956 285592
rect 121696 285552 124956 285580
rect 121696 285540 121702 285552
rect 124950 285540 124956 285552
rect 125008 285540 125014 285592
rect 121546 284316 121552 284368
rect 121604 284356 121610 284368
rect 250438 284356 250444 284368
rect 121604 284328 250444 284356
rect 121604 284316 121610 284328
rect 250438 284316 250444 284328
rect 250496 284316 250502 284368
rect 121638 284180 121644 284232
rect 121696 284220 121702 284232
rect 124858 284220 124864 284232
rect 121696 284192 124864 284220
rect 121696 284180 121702 284192
rect 124858 284180 124864 284192
rect 124916 284180 124922 284232
rect 57790 282888 57796 282940
rect 57848 282928 57854 282940
rect 67634 282928 67640 282940
rect 57848 282900 67640 282928
rect 57848 282888 57854 282900
rect 67634 282888 67640 282900
rect 67692 282888 67698 282940
rect 121454 282888 121460 282940
rect 121512 282928 121518 282940
rect 345014 282928 345020 282940
rect 121512 282900 345020 282928
rect 121512 282888 121518 282900
rect 345014 282888 345020 282900
rect 345072 282888 345078 282940
rect 121454 281596 121460 281648
rect 121512 281636 121518 281648
rect 195238 281636 195244 281648
rect 121512 281608 195244 281636
rect 121512 281596 121518 281608
rect 195238 281596 195244 281608
rect 195296 281596 195302 281648
rect 121638 281528 121644 281580
rect 121696 281568 121702 281580
rect 242158 281568 242164 281580
rect 121696 281540 242164 281568
rect 121696 281528 121702 281540
rect 242158 281528 242164 281540
rect 242216 281528 242222 281580
rect 121454 280236 121460 280288
rect 121512 280276 121518 280288
rect 262214 280276 262220 280288
rect 121512 280248 262220 280276
rect 121512 280236 121518 280248
rect 262214 280236 262220 280248
rect 262272 280236 262278 280288
rect 63402 280168 63408 280220
rect 63460 280208 63466 280220
rect 67634 280208 67640 280220
rect 63460 280180 67640 280208
rect 63460 280168 63466 280180
rect 67634 280168 67640 280180
rect 67692 280168 67698 280220
rect 121638 280168 121644 280220
rect 121696 280208 121702 280220
rect 321554 280208 321560 280220
rect 121696 280180 321560 280208
rect 121696 280168 121702 280180
rect 321554 280168 321560 280180
rect 321612 280168 321618 280220
rect 66162 280100 66168 280152
rect 66220 280140 66226 280152
rect 67726 280140 67732 280152
rect 66220 280112 67732 280140
rect 66220 280100 66226 280112
rect 67726 280100 67732 280112
rect 67784 280100 67790 280152
rect 121454 278808 121460 278860
rect 121512 278848 121518 278860
rect 231118 278848 231124 278860
rect 121512 278820 231124 278848
rect 121512 278808 121518 278820
rect 231118 278808 231124 278820
rect 231176 278808 231182 278860
rect 51718 278740 51724 278792
rect 51776 278780 51782 278792
rect 67634 278780 67640 278792
rect 51776 278752 67640 278780
rect 51776 278740 51782 278752
rect 67634 278740 67640 278752
rect 67692 278740 67698 278792
rect 121638 278740 121644 278792
rect 121696 278780 121702 278792
rect 313918 278780 313924 278792
rect 121696 278752 313924 278780
rect 121696 278740 121702 278752
rect 313918 278740 313924 278752
rect 313976 278740 313982 278792
rect 56410 277448 56416 277500
rect 56468 277488 56474 277500
rect 67634 277488 67640 277500
rect 56468 277460 67640 277488
rect 56468 277448 56474 277460
rect 67634 277448 67640 277460
rect 67692 277448 67698 277500
rect 121638 277448 121644 277500
rect 121696 277488 121702 277500
rect 328454 277488 328460 277500
rect 121696 277460 328460 277488
rect 121696 277448 121702 277460
rect 328454 277448 328460 277460
rect 328512 277448 328518 277500
rect 54938 277380 54944 277432
rect 54996 277420 55002 277432
rect 67726 277420 67732 277432
rect 54996 277392 67732 277420
rect 54996 277380 55002 277392
rect 67726 277380 67732 277392
rect 67784 277380 67790 277432
rect 121454 277380 121460 277432
rect 121512 277420 121518 277432
rect 346486 277420 346492 277432
rect 121512 277392 346492 277420
rect 121512 277380 121518 277392
rect 346486 277380 346492 277392
rect 346544 277380 346550 277432
rect 65886 276088 65892 276140
rect 65944 276128 65950 276140
rect 68002 276128 68008 276140
rect 65944 276100 68008 276128
rect 65944 276088 65950 276100
rect 68002 276088 68008 276100
rect 68060 276088 68066 276140
rect 55030 276020 55036 276072
rect 55088 276060 55094 276072
rect 67634 276060 67640 276072
rect 55088 276032 67640 276060
rect 55088 276020 55094 276032
rect 67634 276020 67640 276032
rect 67692 276020 67698 276072
rect 121454 276020 121460 276072
rect 121512 276060 121518 276072
rect 144178 276060 144184 276072
rect 121512 276032 144184 276060
rect 121512 276020 121518 276032
rect 144178 276020 144184 276032
rect 144236 276020 144242 276072
rect 122282 275272 122288 275324
rect 122340 275312 122346 275324
rect 393958 275312 393964 275324
rect 122340 275284 393964 275312
rect 122340 275272 122346 275284
rect 393958 275272 393964 275284
rect 394016 275272 394022 275324
rect 57698 274660 57704 274712
rect 57756 274700 57762 274712
rect 67634 274700 67640 274712
rect 57756 274672 67640 274700
rect 57756 274660 57762 274672
rect 67634 274660 67640 274672
rect 67692 274660 67698 274712
rect 121454 274660 121460 274712
rect 121512 274700 121518 274712
rect 255498 274700 255504 274712
rect 121512 274672 255504 274700
rect 121512 274660 121518 274672
rect 255498 274660 255504 274672
rect 255556 274660 255562 274712
rect 17218 274592 17224 274644
rect 17276 274632 17282 274644
rect 67726 274632 67732 274644
rect 17276 274604 67732 274632
rect 17276 274592 17282 274604
rect 67726 274592 67732 274604
rect 67784 274592 67790 274644
rect 121454 274252 121460 274304
rect 121512 274292 121518 274304
rect 123662 274292 123668 274304
rect 121512 274264 123668 274292
rect 121512 274252 121518 274264
rect 123662 274252 123668 274264
rect 123720 274252 123726 274304
rect 66070 273232 66076 273284
rect 66128 273272 66134 273284
rect 68002 273272 68008 273284
rect 66128 273244 68008 273272
rect 66128 273232 66134 273244
rect 68002 273232 68008 273244
rect 68060 273232 68066 273284
rect 121454 273232 121460 273284
rect 121512 273272 121518 273284
rect 228358 273272 228364 273284
rect 121512 273244 228364 273272
rect 121512 273232 121518 273244
rect 228358 273232 228364 273244
rect 228416 273232 228422 273284
rect 61930 271940 61936 271992
rect 61988 271980 61994 271992
rect 67634 271980 67640 271992
rect 61988 271952 67640 271980
rect 61988 271940 61994 271952
rect 67634 271940 67640 271952
rect 67692 271940 67698 271992
rect 60550 271872 60556 271924
rect 60608 271912 60614 271924
rect 67726 271912 67732 271924
rect 60608 271884 67732 271912
rect 60608 271872 60614 271884
rect 67726 271872 67732 271884
rect 67784 271872 67790 271924
rect 130470 271872 130476 271924
rect 130528 271912 130534 271924
rect 580166 271912 580172 271924
rect 130528 271884 580172 271912
rect 130528 271872 130534 271884
rect 580166 271872 580172 271884
rect 580224 271872 580230 271924
rect 121638 271124 121644 271176
rect 121696 271164 121702 271176
rect 329926 271164 329932 271176
rect 121696 271136 329932 271164
rect 121696 271124 121702 271136
rect 329926 271124 329932 271136
rect 329984 271124 329990 271176
rect 49602 270512 49608 270564
rect 49660 270552 49666 270564
rect 67634 270552 67640 270564
rect 49660 270524 67640 270552
rect 49660 270512 49666 270524
rect 67634 270512 67640 270524
rect 67692 270512 67698 270564
rect 6914 269764 6920 269816
rect 6972 269804 6978 269816
rect 63494 269804 63500 269816
rect 6972 269776 63500 269804
rect 6972 269764 6978 269776
rect 63494 269764 63500 269776
rect 63552 269764 63558 269816
rect 59170 269084 59176 269136
rect 59228 269124 59234 269136
rect 67634 269124 67640 269136
rect 59228 269096 67640 269124
rect 59228 269084 59234 269096
rect 67634 269084 67640 269096
rect 67692 269084 67698 269136
rect 121454 269084 121460 269136
rect 121512 269124 121518 269136
rect 180058 269124 180064 269136
rect 121512 269096 180064 269124
rect 121512 269084 121518 269096
rect 180058 269084 180064 269096
rect 180116 269084 180122 269136
rect 121546 268336 121552 268388
rect 121604 268376 121610 268388
rect 252646 268376 252652 268388
rect 121604 268348 252652 268376
rect 121604 268336 121610 268348
rect 252646 268336 252652 268348
rect 252704 268336 252710 268388
rect 32398 267724 32404 267776
rect 32456 267764 32462 267776
rect 67634 267764 67640 267776
rect 32456 267736 67640 267764
rect 32456 267724 32462 267736
rect 67634 267724 67640 267736
rect 67692 267724 67698 267776
rect 121454 267724 121460 267776
rect 121512 267764 121518 267776
rect 284938 267764 284944 267776
rect 121512 267736 284944 267764
rect 121512 267724 121518 267736
rect 284938 267724 284944 267736
rect 284996 267724 285002 267776
rect 29638 267656 29644 267708
rect 29696 267696 29702 267708
rect 67726 267696 67732 267708
rect 29696 267668 67732 267696
rect 29696 267656 29702 267668
rect 67726 267656 67732 267668
rect 67784 267656 67790 267708
rect 63494 267588 63500 267640
rect 63552 267628 63558 267640
rect 67634 267628 67640 267640
rect 63552 267600 67640 267628
rect 63552 267588 63558 267600
rect 67634 267588 67640 267600
rect 67692 267588 67698 267640
rect 121638 266976 121644 267028
rect 121696 267016 121702 267028
rect 126330 267016 126336 267028
rect 121696 266988 126336 267016
rect 121696 266976 121702 266988
rect 126330 266976 126336 266988
rect 126388 266976 126394 267028
rect 121454 266432 121460 266484
rect 121512 266472 121518 266484
rect 276658 266472 276664 266484
rect 121512 266444 276664 266472
rect 121512 266432 121518 266444
rect 276658 266432 276664 266444
rect 276716 266432 276722 266484
rect 121546 266364 121552 266416
rect 121604 266404 121610 266416
rect 343726 266404 343732 266416
rect 121604 266376 343732 266404
rect 121604 266364 121610 266376
rect 343726 266364 343732 266376
rect 343784 266364 343790 266416
rect 21358 266296 21364 266348
rect 21416 266336 21422 266348
rect 67726 266336 67732 266348
rect 21416 266308 67732 266336
rect 21416 266296 21422 266308
rect 67726 266296 67732 266308
rect 67784 266296 67790 266348
rect 121454 265004 121460 265056
rect 121512 265044 121518 265056
rect 309778 265044 309784 265056
rect 121512 265016 309784 265044
rect 121512 265004 121518 265016
rect 309778 265004 309784 265016
rect 309836 265004 309842 265056
rect 53650 264936 53656 264988
rect 53708 264976 53714 264988
rect 67634 264976 67640 264988
rect 53708 264948 67640 264976
rect 53708 264936 53714 264948
rect 67634 264936 67640 264948
rect 67692 264936 67698 264988
rect 121546 264936 121552 264988
rect 121604 264976 121610 264988
rect 339586 264976 339592 264988
rect 121604 264948 339592 264976
rect 121604 264936 121610 264948
rect 339586 264936 339592 264948
rect 339644 264936 339650 264988
rect 59262 263644 59268 263696
rect 59320 263684 59326 263696
rect 67634 263684 67640 263696
rect 59320 263656 67640 263684
rect 59320 263644 59326 263656
rect 67634 263644 67640 263656
rect 67692 263644 67698 263696
rect 17218 263576 17224 263628
rect 17276 263616 17282 263628
rect 67726 263616 67732 263628
rect 17276 263588 67732 263616
rect 17276 263576 17282 263588
rect 67726 263576 67732 263588
rect 67784 263576 67790 263628
rect 121546 263576 121552 263628
rect 121604 263616 121610 263628
rect 253934 263616 253940 263628
rect 121604 263588 253940 263616
rect 121604 263576 121610 263588
rect 253934 263576 253940 263588
rect 253992 263576 253998 263628
rect 18598 263508 18604 263560
rect 18656 263548 18662 263560
rect 67634 263548 67640 263560
rect 18656 263520 67640 263548
rect 18656 263508 18662 263520
rect 67634 263508 67640 263520
rect 67692 263508 67698 263560
rect 121454 263508 121460 263560
rect 121512 263548 121518 263560
rect 125594 263548 125600 263560
rect 121512 263520 125600 263548
rect 121512 263508 121518 263520
rect 125594 263508 125600 263520
rect 125652 263508 125658 263560
rect 144178 262828 144184 262880
rect 144236 262868 144242 262880
rect 580350 262868 580356 262880
rect 144236 262840 580356 262868
rect 144236 262828 144242 262840
rect 580350 262828 580356 262840
rect 580408 262828 580414 262880
rect 60458 262216 60464 262268
rect 60516 262256 60522 262268
rect 67634 262256 67640 262268
rect 60516 262228 67640 262256
rect 60516 262216 60522 262228
rect 67634 262216 67640 262228
rect 67692 262216 67698 262268
rect 121454 262216 121460 262268
rect 121512 262256 121518 262268
rect 340874 262256 340880 262268
rect 121512 262228 340880 262256
rect 121512 262216 121518 262228
rect 340874 262216 340880 262228
rect 340932 262216 340938 262268
rect 119798 261468 119804 261520
rect 119856 261508 119862 261520
rect 324590 261508 324596 261520
rect 119856 261480 324596 261508
rect 119856 261468 119862 261480
rect 324590 261468 324596 261480
rect 324648 261468 324654 261520
rect 65978 260924 65984 260976
rect 66036 260964 66042 260976
rect 67634 260964 67640 260976
rect 66036 260936 67640 260964
rect 66036 260924 66042 260936
rect 67634 260924 67640 260936
rect 67692 260924 67698 260976
rect 61838 260856 61844 260908
rect 61896 260896 61902 260908
rect 67726 260896 67732 260908
rect 61896 260868 67732 260896
rect 61896 260856 61902 260868
rect 67726 260856 67732 260868
rect 67784 260856 67790 260908
rect 121454 260856 121460 260908
rect 121512 260896 121518 260908
rect 343634 260896 343640 260908
rect 121512 260868 343640 260896
rect 121512 260856 121518 260868
rect 343634 260856 343640 260868
rect 343692 260856 343698 260908
rect 39298 260788 39304 260840
rect 39356 260828 39362 260840
rect 67634 260828 67640 260840
rect 39356 260800 67640 260828
rect 39356 260788 39362 260800
rect 67634 260788 67640 260800
rect 67692 260788 67698 260840
rect 56502 259428 56508 259480
rect 56560 259468 56566 259480
rect 67634 259468 67640 259480
rect 56560 259440 67640 259468
rect 56560 259428 56566 259440
rect 67634 259428 67640 259440
rect 67692 259428 67698 259480
rect 121454 259428 121460 259480
rect 121512 259468 121518 259480
rect 246298 259468 246304 259480
rect 121512 259440 246304 259468
rect 121512 259428 121518 259440
rect 246298 259428 246304 259440
rect 246356 259428 246362 259480
rect 121546 259360 121552 259412
rect 121604 259400 121610 259412
rect 151078 259400 151084 259412
rect 121604 259372 151084 259400
rect 121604 259360 121610 259372
rect 151078 259360 151084 259372
rect 151136 259360 151142 259412
rect 342898 259360 342904 259412
rect 342956 259400 342962 259412
rect 579798 259400 579804 259412
rect 342956 259372 579804 259400
rect 342956 259360 342962 259372
rect 579798 259360 579804 259372
rect 579856 259360 579862 259412
rect 64782 258136 64788 258188
rect 64840 258176 64846 258188
rect 67634 258176 67640 258188
rect 64840 258148 67640 258176
rect 64840 258136 64846 258148
rect 67634 258136 67640 258148
rect 67692 258136 67698 258188
rect 57514 258068 57520 258120
rect 57572 258108 57578 258120
rect 67726 258108 67732 258120
rect 57572 258080 67732 258108
rect 57572 258068 57578 258080
rect 67726 258068 67732 258080
rect 67784 258068 67790 258120
rect 121454 258068 121460 258120
rect 121512 258108 121518 258120
rect 331214 258108 331220 258120
rect 121512 258080 331220 258108
rect 121512 258068 121518 258080
rect 331214 258068 331220 258080
rect 331272 258068 331278 258120
rect 121454 257864 121460 257916
rect 121512 257904 121518 257916
rect 125042 257904 125048 257916
rect 121512 257876 125048 257904
rect 121512 257864 121518 257876
rect 125042 257864 125048 257876
rect 125100 257864 125106 257916
rect 50982 257320 50988 257372
rect 51040 257360 51046 257372
rect 68278 257360 68284 257372
rect 51040 257332 68284 257360
rect 51040 257320 51046 257332
rect 68278 257320 68284 257332
rect 68336 257320 68342 257372
rect 124858 257320 124864 257372
rect 124916 257360 124922 257372
rect 582374 257360 582380 257372
rect 124916 257332 582380 257360
rect 124916 257320 124922 257332
rect 582374 257320 582380 257332
rect 582432 257320 582438 257372
rect 14458 256708 14464 256760
rect 14516 256748 14522 256760
rect 67634 256748 67640 256760
rect 14516 256720 67640 256748
rect 14516 256708 14522 256720
rect 67634 256708 67640 256720
rect 67692 256708 67698 256760
rect 121546 256708 121552 256760
rect 121604 256748 121610 256760
rect 232498 256748 232504 256760
rect 121604 256720 232504 256748
rect 121604 256708 121610 256720
rect 232498 256708 232504 256720
rect 232556 256708 232562 256760
rect 121638 256640 121644 256692
rect 121696 256680 121702 256692
rect 130378 256680 130384 256692
rect 121696 256652 130384 256680
rect 121696 256640 121702 256652
rect 130378 256640 130384 256652
rect 130436 256640 130442 256692
rect 121454 256572 121460 256624
rect 121512 256612 121518 256624
rect 129090 256612 129096 256624
rect 121512 256584 129096 256612
rect 121512 256572 121518 256584
rect 129090 256572 129096 256584
rect 129148 256572 129154 256624
rect 64598 255348 64604 255400
rect 64656 255388 64662 255400
rect 67634 255388 67640 255400
rect 64656 255360 67640 255388
rect 64656 255348 64662 255360
rect 67634 255348 67640 255360
rect 67692 255348 67698 255400
rect 60642 255280 60648 255332
rect 60700 255320 60706 255332
rect 67726 255320 67732 255332
rect 60700 255292 67732 255320
rect 60700 255280 60706 255292
rect 67726 255280 67732 255292
rect 67784 255280 67790 255332
rect 57882 255212 57888 255264
rect 57940 255252 57946 255264
rect 67634 255252 67640 255264
rect 57940 255224 67640 255252
rect 57940 255212 57946 255224
rect 67634 255212 67640 255224
rect 67692 255212 67698 255264
rect 121454 253988 121460 254040
rect 121512 254028 121518 254040
rect 273254 254028 273260 254040
rect 121512 254000 273260 254028
rect 121512 253988 121518 254000
rect 273254 253988 273260 254000
rect 273312 253988 273318 254040
rect 3142 253920 3148 253972
rect 3200 253960 3206 253972
rect 18598 253960 18604 253972
rect 3200 253932 18604 253960
rect 3200 253920 3206 253932
rect 18598 253920 18604 253932
rect 18656 253920 18662 253972
rect 121546 253920 121552 253972
rect 121604 253960 121610 253972
rect 327074 253960 327080 253972
rect 121604 253932 327080 253960
rect 121604 253920 121610 253932
rect 327074 253920 327080 253932
rect 327132 253920 327138 253972
rect 64690 252628 64696 252680
rect 64748 252668 64754 252680
rect 67634 252668 67640 252680
rect 64748 252640 67640 252668
rect 64748 252628 64754 252640
rect 67634 252628 67640 252640
rect 67692 252628 67698 252680
rect 22738 252560 22744 252612
rect 22796 252600 22802 252612
rect 67726 252600 67732 252612
rect 22796 252572 67732 252600
rect 22796 252560 22802 252572
rect 67726 252560 67732 252572
rect 67784 252560 67790 252612
rect 121546 252560 121552 252612
rect 121604 252600 121610 252612
rect 316678 252600 316684 252612
rect 121604 252572 316684 252600
rect 121604 252560 121610 252572
rect 316678 252560 316684 252572
rect 316736 252560 316742 252612
rect 121454 252492 121460 252544
rect 121512 252532 121518 252544
rect 126238 252532 126244 252544
rect 121512 252504 126244 252532
rect 121512 252492 121518 252504
rect 126238 252492 126244 252504
rect 126296 252492 126302 252544
rect 63310 251200 63316 251252
rect 63368 251240 63374 251252
rect 67634 251240 67640 251252
rect 63368 251212 67640 251240
rect 63368 251200 63374 251212
rect 67634 251200 67640 251212
rect 67692 251200 67698 251252
rect 121454 250452 121460 250504
rect 121512 250492 121518 250504
rect 327166 250492 327172 250504
rect 121512 250464 327172 250492
rect 121512 250452 121518 250464
rect 327166 250452 327172 250464
rect 327224 250452 327230 250504
rect 60366 249840 60372 249892
rect 60424 249880 60430 249892
rect 67634 249880 67640 249892
rect 60424 249852 67640 249880
rect 60424 249840 60430 249852
rect 67634 249840 67640 249852
rect 67692 249840 67698 249892
rect 58986 249772 58992 249824
rect 59044 249812 59050 249824
rect 67726 249812 67732 249824
rect 59044 249784 67732 249812
rect 59044 249772 59050 249784
rect 67726 249772 67732 249784
rect 67784 249772 67790 249824
rect 121546 249772 121552 249824
rect 121604 249812 121610 249824
rect 209038 249812 209044 249824
rect 121604 249784 209044 249812
rect 121604 249772 121610 249784
rect 209038 249772 209044 249784
rect 209096 249772 209102 249824
rect 62022 249704 62028 249756
rect 62080 249744 62086 249756
rect 67634 249744 67640 249756
rect 62080 249716 67640 249744
rect 62080 249704 62086 249716
rect 67634 249704 67640 249716
rect 67692 249704 67698 249756
rect 121454 249704 121460 249756
rect 121512 249744 121518 249756
rect 141418 249744 141424 249756
rect 121512 249716 141424 249744
rect 121512 249704 121518 249716
rect 141418 249704 141424 249716
rect 141476 249704 141482 249756
rect 67542 249636 67548 249688
rect 67600 249676 67606 249688
rect 68370 249676 68376 249688
rect 67600 249648 68376 249676
rect 67600 249636 67606 249648
rect 68370 249636 68376 249648
rect 68428 249636 68434 249688
rect 57606 248412 57612 248464
rect 57664 248452 57670 248464
rect 67634 248452 67640 248464
rect 57664 248424 67640 248452
rect 57664 248412 57670 248424
rect 67634 248412 67640 248424
rect 67692 248412 67698 248464
rect 121454 248412 121460 248464
rect 121512 248452 121518 248464
rect 353294 248452 353300 248464
rect 121512 248424 353300 248452
rect 121512 248412 121518 248424
rect 353294 248412 353300 248424
rect 353352 248412 353358 248464
rect 62022 247120 62028 247172
rect 62080 247160 62086 247172
rect 67634 247160 67640 247172
rect 62080 247132 67640 247160
rect 62080 247120 62086 247132
rect 67634 247120 67640 247132
rect 67692 247120 67698 247172
rect 61746 247052 61752 247104
rect 61804 247092 61810 247104
rect 67726 247092 67732 247104
rect 61804 247064 67732 247092
rect 61804 247052 61810 247064
rect 67726 247052 67732 247064
rect 67784 247052 67790 247104
rect 121454 247052 121460 247104
rect 121512 247092 121518 247104
rect 263594 247092 263600 247104
rect 121512 247064 263600 247092
rect 121512 247052 121518 247064
rect 263594 247052 263600 247064
rect 263652 247052 263658 247104
rect 53742 246984 53748 247036
rect 53800 247024 53806 247036
rect 67634 247024 67640 247036
rect 53800 246996 67640 247024
rect 53800 246984 53806 246996
rect 67634 246984 67640 246996
rect 67692 246984 67698 247036
rect 64506 245624 64512 245676
rect 64564 245664 64570 245676
rect 67726 245664 67732 245676
rect 64564 245636 67732 245664
rect 64564 245624 64570 245636
rect 67726 245624 67732 245636
rect 67784 245624 67790 245676
rect 121546 245624 121552 245676
rect 121604 245664 121610 245676
rect 266446 245664 266452 245676
rect 121604 245636 266452 245664
rect 121604 245624 121610 245636
rect 266446 245624 266452 245636
rect 266504 245624 266510 245676
rect 33778 245556 33784 245608
rect 33836 245596 33842 245608
rect 67634 245596 67640 245608
rect 33836 245568 67640 245596
rect 33836 245556 33842 245568
rect 67634 245556 67640 245568
rect 67692 245556 67698 245608
rect 121454 245556 121460 245608
rect 121512 245596 121518 245608
rect 128998 245596 129004 245608
rect 121512 245568 129004 245596
rect 121512 245556 121518 245568
rect 128998 245556 129004 245568
rect 129056 245556 129062 245608
rect 121546 244332 121552 244384
rect 121604 244372 121610 244384
rect 289078 244372 289084 244384
rect 121604 244344 289084 244372
rect 121604 244332 121610 244344
rect 289078 244332 289084 244344
rect 289136 244332 289142 244384
rect 63218 244264 63224 244316
rect 63276 244304 63282 244316
rect 67634 244304 67640 244316
rect 63276 244276 67640 244304
rect 63276 244264 63282 244276
rect 67634 244264 67640 244276
rect 67692 244264 67698 244316
rect 128354 244264 128360 244316
rect 128412 244304 128418 244316
rect 579890 244304 579896 244316
rect 128412 244276 579896 244304
rect 128412 244264 128418 244276
rect 579890 244264 579896 244276
rect 579948 244264 579954 244316
rect 4798 244196 4804 244248
rect 4856 244236 4862 244248
rect 67726 244236 67732 244248
rect 4856 244208 67732 244236
rect 4856 244196 4862 244208
rect 67726 244196 67732 244208
rect 67784 244196 67790 244248
rect 121454 244196 121460 244248
rect 121512 244236 121518 244248
rect 134518 244236 134524 244248
rect 121512 244208 134524 244236
rect 121512 244196 121518 244208
rect 134518 244196 134524 244208
rect 134576 244196 134582 244248
rect 122098 243516 122104 243568
rect 122156 243556 122162 243568
rect 238018 243556 238024 243568
rect 122156 243528 238024 243556
rect 122156 243516 122162 243528
rect 238018 243516 238024 243528
rect 238076 243516 238082 243568
rect 121546 242836 121552 242888
rect 121604 242876 121610 242888
rect 133138 242876 133144 242888
rect 121604 242848 133144 242876
rect 121604 242836 121610 242848
rect 133138 242836 133144 242848
rect 133196 242836 133202 242888
rect 121454 242768 121460 242820
rect 121512 242808 121518 242820
rect 128354 242808 128360 242820
rect 121512 242780 128360 242808
rect 121512 242768 121518 242780
rect 128354 242768 128360 242780
rect 128412 242768 128418 242820
rect 160738 242224 160744 242276
rect 160796 242264 160802 242276
rect 318058 242264 318064 242276
rect 160796 242236 318064 242264
rect 160796 242224 160802 242236
rect 318058 242224 318064 242236
rect 318116 242224 318122 242276
rect 121638 242156 121644 242208
rect 121696 242196 121702 242208
rect 327258 242196 327264 242208
rect 121696 242168 327264 242196
rect 121696 242156 121702 242168
rect 327258 242156 327264 242168
rect 327316 242156 327322 242208
rect 63126 241476 63132 241528
rect 63184 241516 63190 241528
rect 67634 241516 67640 241528
rect 63184 241488 67640 241516
rect 63184 241476 63190 241488
rect 67634 241476 67640 241488
rect 67692 241476 67698 241528
rect 121454 240184 121460 240236
rect 121512 240224 121518 240236
rect 222838 240224 222844 240236
rect 121512 240196 222844 240224
rect 121512 240184 121518 240196
rect 222838 240184 222844 240196
rect 222896 240184 222902 240236
rect 3050 240116 3056 240168
rect 3108 240156 3114 240168
rect 15194 240156 15200 240168
rect 3108 240128 15200 240156
rect 3108 240116 3114 240128
rect 15194 240116 15200 240128
rect 15252 240116 15258 240168
rect 121546 240116 121552 240168
rect 121604 240156 121610 240168
rect 330018 240156 330024 240168
rect 121604 240128 330024 240156
rect 121604 240116 121610 240128
rect 330018 240116 330024 240128
rect 330076 240116 330082 240168
rect 118326 239912 118332 239964
rect 118384 239952 118390 239964
rect 123478 239952 123484 239964
rect 118384 239924 123484 239952
rect 118384 239912 118390 239924
rect 123478 239912 123484 239924
rect 123536 239912 123542 239964
rect 73154 239776 73160 239828
rect 73212 239816 73218 239828
rect 73878 239816 73884 239828
rect 73212 239788 73884 239816
rect 73212 239776 73218 239788
rect 73878 239776 73884 239788
rect 73936 239776 73942 239828
rect 75914 239776 75920 239828
rect 75972 239816 75978 239828
rect 77098 239816 77104 239828
rect 75972 239788 77104 239816
rect 75972 239776 75978 239788
rect 77098 239776 77104 239788
rect 77156 239776 77162 239828
rect 77294 239776 77300 239828
rect 77352 239816 77358 239828
rect 78386 239816 78392 239828
rect 77352 239788 78392 239816
rect 77352 239776 77358 239788
rect 78386 239776 78392 239788
rect 78444 239776 78450 239828
rect 78674 239776 78680 239828
rect 78732 239816 78738 239828
rect 79674 239816 79680 239828
rect 78732 239788 79680 239816
rect 78732 239776 78738 239788
rect 79674 239776 79680 239788
rect 79732 239776 79738 239828
rect 82814 239776 82820 239828
rect 82872 239816 82878 239828
rect 83538 239816 83544 239828
rect 82872 239788 83544 239816
rect 82872 239776 82878 239788
rect 83538 239776 83544 239788
rect 83596 239776 83602 239828
rect 86954 239776 86960 239828
rect 87012 239816 87018 239828
rect 88046 239816 88052 239828
rect 87012 239788 88052 239816
rect 87012 239776 87018 239788
rect 88046 239776 88052 239788
rect 88104 239776 88110 239828
rect 89714 239776 89720 239828
rect 89772 239816 89778 239828
rect 90622 239816 90628 239828
rect 89772 239788 90628 239816
rect 89772 239776 89778 239788
rect 90622 239776 90628 239788
rect 90680 239776 90686 239828
rect 92474 239776 92480 239828
rect 92532 239816 92538 239828
rect 93198 239816 93204 239828
rect 92532 239788 93204 239816
rect 92532 239776 92538 239788
rect 93198 239776 93204 239788
rect 93256 239776 93262 239828
rect 104894 239776 104900 239828
rect 104952 239816 104958 239828
rect 106078 239816 106084 239828
rect 104952 239788 106084 239816
rect 104952 239776 104958 239788
rect 106078 239776 106084 239788
rect 106136 239776 106142 239828
rect 114554 239776 114560 239828
rect 114612 239816 114618 239828
rect 115738 239816 115744 239828
rect 114612 239788 115744 239816
rect 114612 239776 114618 239788
rect 115738 239776 115744 239788
rect 115796 239776 115802 239828
rect 64690 239504 64696 239556
rect 64748 239544 64754 239556
rect 72418 239544 72424 239556
rect 64748 239516 72424 239544
rect 64748 239504 64754 239516
rect 72418 239504 72424 239516
rect 72476 239504 72482 239556
rect 63310 239436 63316 239488
rect 63368 239476 63374 239488
rect 98638 239476 98644 239488
rect 63368 239448 98644 239476
rect 63368 239436 63374 239448
rect 98638 239436 98644 239448
rect 98696 239436 98702 239488
rect 3602 239368 3608 239420
rect 3660 239408 3666 239420
rect 63494 239408 63500 239420
rect 3660 239380 63500 239408
rect 3660 239368 3666 239380
rect 63494 239368 63500 239380
rect 63552 239368 63558 239420
rect 69658 239368 69664 239420
rect 69716 239408 69722 239420
rect 312538 239408 312544 239420
rect 69716 239380 312544 239408
rect 69716 239368 69722 239380
rect 312538 239368 312544 239380
rect 312596 239368 312602 239420
rect 84286 239300 84292 239352
rect 84344 239340 84350 239352
rect 85482 239340 85488 239352
rect 84344 239312 85488 239340
rect 84344 239300 84350 239312
rect 85482 239300 85488 239312
rect 85540 239300 85546 239352
rect 106734 238756 106740 238808
rect 106792 238796 106798 238808
rect 266354 238796 266360 238808
rect 106792 238768 266360 238796
rect 106792 238756 106798 238768
rect 266354 238756 266360 238768
rect 266412 238756 266418 238808
rect 15194 238688 15200 238740
rect 15252 238728 15258 238740
rect 103514 238728 103520 238740
rect 15252 238700 103520 238728
rect 15252 238688 15258 238700
rect 103514 238688 103520 238700
rect 103572 238688 103578 238740
rect 113818 238688 113824 238740
rect 113876 238728 113882 238740
rect 305638 238728 305644 238740
rect 113876 238700 305644 238728
rect 113876 238688 113882 238700
rect 305638 238688 305644 238700
rect 305696 238688 305702 238740
rect 40034 238620 40040 238672
rect 40092 238660 40098 238672
rect 95786 238660 95792 238672
rect 40092 238632 95792 238660
rect 40092 238620 40098 238632
rect 95786 238620 95792 238632
rect 95844 238620 95850 238672
rect 117038 238620 117044 238672
rect 117096 238660 117102 238672
rect 124858 238660 124864 238672
rect 117096 238632 124864 238660
rect 117096 238620 117102 238632
rect 124858 238620 124864 238632
rect 124916 238620 124922 238672
rect 52362 238552 52368 238604
rect 52420 238592 52426 238604
rect 75822 238592 75828 238604
rect 52420 238564 75828 238592
rect 52420 238552 52426 238564
rect 75822 238552 75828 238564
rect 75880 238552 75886 238604
rect 91278 238552 91284 238604
rect 91336 238592 91342 238604
rect 130470 238592 130476 238604
rect 91336 238564 130476 238592
rect 91336 238552 91342 238564
rect 130470 238552 130476 238564
rect 130528 238552 130534 238604
rect 63494 238484 63500 238536
rect 63552 238524 63558 238536
rect 86770 238524 86776 238536
rect 63552 238496 86776 238524
rect 63552 238484 63558 238496
rect 86770 238484 86776 238496
rect 86828 238484 86834 238536
rect 115106 238484 115112 238536
rect 115164 238524 115170 238536
rect 123570 238524 123576 238536
rect 115164 238496 123576 238524
rect 115164 238484 115170 238496
rect 123570 238484 123576 238496
rect 123628 238484 123634 238536
rect 102870 238212 102876 238264
rect 102928 238252 102934 238264
rect 106918 238252 106924 238264
rect 102928 238224 106924 238252
rect 102928 238212 102934 238224
rect 106918 238212 106924 238224
rect 106976 238212 106982 238264
rect 81618 238144 81624 238196
rect 81676 238184 81682 238196
rect 114830 238184 114836 238196
rect 81676 238156 114836 238184
rect 81676 238144 81682 238156
rect 114830 238144 114836 238156
rect 114888 238144 114894 238196
rect 72602 238076 72608 238128
rect 72660 238116 72666 238128
rect 91094 238116 91100 238128
rect 72660 238088 91100 238116
rect 72660 238076 72666 238088
rect 91094 238076 91100 238088
rect 91152 238076 91158 238128
rect 105446 238076 105452 238128
rect 105504 238116 105510 238128
rect 196618 238116 196624 238128
rect 105504 238088 196624 238116
rect 105504 238076 105510 238088
rect 196618 238076 196624 238088
rect 196676 238076 196682 238128
rect 71314 238008 71320 238060
rect 71372 238048 71378 238060
rect 79318 238048 79324 238060
rect 71372 238020 79324 238048
rect 71372 238008 71378 238020
rect 79318 238008 79324 238020
rect 79376 238008 79382 238060
rect 86126 238008 86132 238060
rect 86184 238048 86190 238060
rect 582374 238048 582380 238060
rect 86184 238020 582380 238048
rect 86184 238008 86190 238020
rect 582374 238008 582380 238020
rect 582432 238008 582438 238060
rect 35158 237328 35164 237380
rect 35216 237368 35222 237380
rect 82262 237368 82268 237380
rect 35216 237340 82268 237368
rect 35216 237328 35222 237340
rect 82262 237328 82268 237340
rect 82320 237328 82326 237380
rect 98362 237328 98368 237380
rect 98420 237368 98426 237380
rect 359458 237368 359464 237380
rect 98420 237340 359464 237368
rect 98420 237328 98426 237340
rect 359458 237328 359464 237340
rect 359516 237328 359522 237380
rect 47578 237260 47584 237312
rect 47636 237300 47642 237312
rect 114462 237300 114468 237312
rect 47636 237272 114468 237300
rect 47636 237260 47642 237272
rect 114462 237260 114468 237272
rect 114520 237260 114526 237312
rect 55122 237192 55128 237244
rect 55180 237232 55186 237244
rect 89346 237232 89352 237244
rect 55180 237204 89352 237232
rect 55180 237192 55186 237204
rect 89346 237192 89352 237204
rect 89404 237192 89410 237244
rect 67358 236648 67364 236700
rect 67416 236688 67422 236700
rect 214650 236688 214656 236700
rect 67416 236660 214656 236688
rect 67416 236648 67422 236660
rect 214650 236648 214656 236660
rect 214708 236648 214714 236700
rect 18598 235900 18604 235952
rect 18656 235940 18662 235952
rect 112530 235940 112536 235952
rect 18656 235912 112536 235940
rect 18656 235900 18662 235912
rect 112530 235900 112536 235912
rect 112588 235900 112594 235952
rect 43438 235832 43444 235884
rect 43496 235872 43502 235884
rect 99006 235872 99012 235884
rect 43496 235844 99012 235872
rect 43496 235832 43502 235844
rect 99006 235832 99012 235844
rect 99064 235832 99070 235884
rect 80330 235288 80336 235340
rect 80388 235328 80394 235340
rect 320818 235328 320824 235340
rect 80388 235300 320824 235328
rect 80388 235288 80394 235300
rect 320818 235288 320824 235300
rect 320876 235288 320882 235340
rect 117682 235220 117688 235272
rect 117740 235260 117746 235272
rect 583110 235260 583116 235272
rect 117740 235232 583116 235260
rect 117740 235220 117746 235232
rect 583110 235220 583116 235232
rect 583168 235220 583174 235272
rect 91922 234540 91928 234592
rect 91980 234580 91986 234592
rect 582650 234580 582656 234592
rect 91980 234552 582656 234580
rect 91980 234540 91986 234552
rect 582650 234540 582656 234552
rect 582708 234540 582714 234592
rect 69014 233928 69020 233980
rect 69072 233968 69078 233980
rect 69750 233968 69756 233980
rect 69072 233940 69756 233968
rect 69072 233928 69078 233940
rect 69750 233928 69756 233940
rect 69808 233928 69814 233980
rect 63218 233860 63224 233912
rect 63276 233900 63282 233912
rect 191190 233900 191196 233912
rect 63276 233872 191196 233900
rect 63276 233860 63282 233872
rect 191190 233860 191196 233872
rect 191248 233860 191254 233912
rect 93854 233724 93860 233776
rect 93912 233764 93918 233776
rect 94038 233764 94044 233776
rect 93912 233736 94044 233764
rect 93912 233724 93918 233736
rect 94038 233724 94044 233736
rect 94096 233724 94102 233776
rect 114830 233180 114836 233232
rect 114888 233220 114894 233232
rect 214558 233220 214564 233232
rect 114888 233192 214564 233220
rect 114888 233180 114894 233192
rect 214558 233180 214564 233192
rect 214616 233180 214622 233232
rect 69198 232500 69204 232552
rect 69256 232540 69262 232552
rect 251174 232540 251180 232552
rect 69256 232512 251180 232540
rect 69256 232500 69262 232512
rect 251174 232500 251180 232512
rect 251232 232500 251238 232552
rect 84102 231820 84108 231872
rect 84160 231860 84166 231872
rect 84838 231860 84844 231872
rect 84160 231832 84844 231860
rect 84160 231820 84166 231832
rect 84838 231820 84844 231832
rect 84896 231820 84902 231872
rect 106826 231752 106832 231804
rect 106884 231792 106890 231804
rect 542354 231792 542360 231804
rect 106884 231764 542360 231792
rect 106884 231752 106890 231764
rect 542354 231752 542360 231764
rect 542412 231752 542418 231804
rect 60366 231208 60372 231260
rect 60424 231248 60430 231260
rect 160738 231248 160744 231260
rect 60424 231220 160744 231248
rect 60424 231208 60430 231220
rect 160738 231208 160744 231220
rect 160796 231208 160802 231260
rect 15838 231140 15844 231192
rect 15896 231180 15902 231192
rect 109862 231180 109868 231192
rect 15896 231152 109868 231180
rect 15896 231140 15902 231152
rect 109862 231140 109868 231152
rect 109920 231140 109926 231192
rect 111794 231140 111800 231192
rect 111852 231180 111858 231192
rect 276014 231180 276020 231192
rect 111852 231152 276020 231180
rect 111852 231140 111858 231152
rect 276014 231140 276020 231152
rect 276072 231140 276078 231192
rect 108574 231072 108580 231124
rect 108632 231112 108638 231124
rect 328546 231112 328552 231124
rect 108632 231084 328552 231112
rect 108632 231072 108638 231084
rect 328546 231072 328552 231084
rect 328604 231072 328610 231124
rect 91094 230392 91100 230444
rect 91152 230432 91158 230444
rect 582558 230432 582564 230444
rect 91152 230404 582564 230432
rect 91152 230392 91158 230404
rect 582558 230392 582564 230404
rect 582616 230392 582622 230444
rect 67266 228420 67272 228472
rect 67324 228460 67330 228472
rect 315298 228460 315304 228472
rect 67324 228432 315304 228460
rect 67324 228420 67330 228432
rect 315298 228420 315304 228432
rect 315356 228420 315362 228472
rect 76006 228352 76012 228404
rect 76064 228392 76070 228404
rect 582558 228392 582564 228404
rect 76064 228364 582564 228392
rect 76064 228352 76070 228364
rect 582558 228352 582564 228364
rect 582616 228352 582622 228404
rect 54938 225564 54944 225616
rect 54996 225604 55002 225616
rect 305638 225604 305644 225616
rect 54996 225576 305644 225604
rect 54996 225564 55002 225576
rect 305638 225564 305644 225576
rect 305696 225564 305702 225616
rect 82906 224272 82912 224324
rect 82964 224312 82970 224324
rect 184198 224312 184204 224324
rect 82964 224284 184204 224312
rect 82964 224272 82970 224284
rect 184198 224272 184204 224284
rect 184256 224272 184262 224324
rect 97626 224204 97632 224256
rect 97684 224244 97690 224256
rect 342346 224244 342352 224256
rect 97684 224216 342352 224244
rect 97684 224204 97690 224216
rect 342346 224204 342352 224216
rect 342404 224204 342410 224256
rect 84286 222844 84292 222896
rect 84344 222884 84350 222896
rect 254118 222884 254124 222896
rect 84344 222856 254124 222884
rect 84344 222844 84350 222856
rect 254118 222844 254124 222856
rect 254176 222844 254182 222896
rect 89806 221484 89812 221536
rect 89864 221524 89870 221536
rect 252738 221524 252744 221536
rect 89864 221496 252744 221524
rect 89864 221484 89870 221496
rect 252738 221484 252744 221496
rect 252796 221484 252802 221536
rect 61838 221416 61844 221468
rect 61896 221456 61902 221468
rect 334066 221456 334072 221468
rect 61896 221428 334072 221456
rect 61896 221416 61902 221428
rect 334066 221416 334072 221428
rect 334124 221416 334130 221468
rect 1302 220192 1308 220244
rect 1360 220232 1366 220244
rect 119798 220232 119804 220244
rect 1360 220204 119804 220232
rect 1360 220192 1366 220204
rect 119798 220192 119804 220204
rect 119856 220192 119862 220244
rect 115934 220124 115940 220176
rect 115992 220164 115998 220176
rect 259730 220164 259736 220176
rect 115992 220136 259736 220164
rect 115992 220124 115998 220136
rect 259730 220124 259736 220136
rect 259788 220124 259794 220176
rect 113358 220056 113364 220108
rect 113416 220096 113422 220108
rect 304258 220096 304264 220108
rect 113416 220068 304264 220096
rect 113416 220056 113422 220068
rect 304258 220056 304264 220068
rect 304316 220056 304322 220108
rect 77386 218696 77392 218748
rect 77444 218736 77450 218748
rect 330110 218736 330116 218748
rect 77444 218708 330116 218736
rect 77444 218696 77450 218708
rect 330110 218696 330116 218708
rect 330168 218696 330174 218748
rect 137278 217404 137284 217456
rect 137336 217444 137342 217456
rect 245010 217444 245016 217456
rect 137336 217416 245016 217444
rect 137336 217404 137342 217416
rect 245010 217404 245016 217416
rect 245068 217404 245074 217456
rect 53650 217336 53656 217388
rect 53708 217376 53714 217388
rect 298738 217376 298744 217388
rect 53708 217348 298744 217376
rect 53708 217336 53714 217348
rect 298738 217336 298744 217348
rect 298796 217336 298802 217388
rect 75914 217268 75920 217320
rect 75972 217308 75978 217320
rect 321646 217308 321652 217320
rect 75972 217280 321652 217308
rect 75972 217268 75978 217280
rect 321646 217268 321652 217280
rect 321704 217268 321710 217320
rect 78766 215976 78772 216028
rect 78824 216016 78830 216028
rect 273346 216016 273352 216028
rect 78824 215988 273352 216016
rect 78824 215976 78830 215988
rect 273346 215976 273352 215988
rect 273404 215976 273410 216028
rect 94038 215908 94044 215960
rect 94096 215948 94102 215960
rect 300118 215948 300124 215960
rect 94096 215920 300124 215948
rect 94096 215908 94102 215920
rect 300118 215908 300124 215920
rect 300176 215908 300182 215960
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 17218 215268 17224 215280
rect 3384 215240 17224 215268
rect 3384 215228 3390 215240
rect 17218 215228 17224 215240
rect 17276 215228 17282 215280
rect 100846 214616 100852 214668
rect 100904 214656 100910 214668
rect 254026 214656 254032 214668
rect 100904 214628 254032 214656
rect 100904 214616 100910 214628
rect 254026 214616 254032 214628
rect 254084 214616 254090 214668
rect 74626 214548 74632 214600
rect 74684 214588 74690 214600
rect 323118 214588 323124 214600
rect 74684 214560 323124 214588
rect 74684 214548 74690 214560
rect 323118 214548 323124 214560
rect 323176 214548 323182 214600
rect 60458 213188 60464 213240
rect 60516 213228 60522 213240
rect 233970 213228 233976 213240
rect 60516 213200 233976 213228
rect 60516 213188 60522 213200
rect 233970 213188 233976 213200
rect 234028 213188 234034 213240
rect 110506 211828 110512 211880
rect 110564 211868 110570 211880
rect 238110 211868 238116 211880
rect 110564 211840 238116 211868
rect 110564 211828 110570 211840
rect 238110 211828 238116 211840
rect 238168 211828 238174 211880
rect 96614 211760 96620 211812
rect 96672 211800 96678 211812
rect 260926 211800 260932 211812
rect 96672 211772 260932 211800
rect 96672 211760 96678 211772
rect 260926 211760 260932 211772
rect 260984 211760 260990 211812
rect 146938 210468 146944 210520
rect 146996 210508 147002 210520
rect 271874 210508 271880 210520
rect 146996 210480 271880 210508
rect 146996 210468 147002 210480
rect 271874 210468 271880 210480
rect 271932 210468 271938 210520
rect 61746 210400 61752 210452
rect 61804 210440 61810 210452
rect 240778 210440 240784 210452
rect 61804 210412 240784 210440
rect 61804 210400 61810 210412
rect 240778 210400 240784 210412
rect 240836 210400 240842 210452
rect 93946 209108 93952 209160
rect 94004 209148 94010 209160
rect 278774 209148 278780 209160
rect 94004 209120 278780 209148
rect 94004 209108 94010 209120
rect 278774 209108 278780 209120
rect 278832 209108 278838 209160
rect 61930 209040 61936 209092
rect 61988 209080 61994 209092
rect 270678 209080 270684 209092
rect 61988 209052 270684 209080
rect 61988 209040 61994 209052
rect 270678 209040 270684 209052
rect 270736 209040 270742 209092
rect 56410 207748 56416 207800
rect 56468 207788 56474 207800
rect 264974 207788 264980 207800
rect 56468 207760 264980 207788
rect 56468 207748 56474 207760
rect 264974 207748 264980 207760
rect 265032 207748 265038 207800
rect 57606 207680 57612 207732
rect 57664 207720 57670 207732
rect 277486 207720 277492 207732
rect 57664 207692 277492 207720
rect 57664 207680 57670 207692
rect 277486 207680 277492 207692
rect 277544 207680 277550 207732
rect 78674 207612 78680 207664
rect 78732 207652 78738 207664
rect 335446 207652 335452 207664
rect 78732 207624 335452 207652
rect 78732 207612 78738 207624
rect 335446 207612 335452 207624
rect 335504 207612 335510 207664
rect 127710 206932 127716 206984
rect 127768 206972 127774 206984
rect 580166 206972 580172 206984
rect 127768 206944 580172 206972
rect 127768 206932 127774 206944
rect 580166 206932 580172 206944
rect 580224 206932 580230 206984
rect 77294 206320 77300 206372
rect 77352 206360 77358 206372
rect 263686 206360 263692 206372
rect 77352 206332 263692 206360
rect 77352 206320 77358 206332
rect 263686 206320 263692 206332
rect 263744 206320 263750 206372
rect 98638 206252 98644 206304
rect 98696 206292 98702 206304
rect 332870 206292 332876 206304
rect 98696 206264 332876 206292
rect 98696 206252 98702 206264
rect 332870 206252 332876 206264
rect 332928 206252 332934 206304
rect 103606 205028 103612 205080
rect 103664 205068 103670 205080
rect 191098 205068 191104 205080
rect 103664 205040 191104 205068
rect 103664 205028 103670 205040
rect 191098 205028 191104 205040
rect 191156 205028 191162 205080
rect 148318 204960 148324 205012
rect 148376 205000 148382 205012
rect 343818 205000 343824 205012
rect 148376 204972 343824 205000
rect 148376 204960 148382 204972
rect 343818 204960 343824 204972
rect 343876 204960 343882 205012
rect 63402 204892 63408 204944
rect 63460 204932 63466 204944
rect 266354 204932 266360 204944
rect 63460 204904 266360 204932
rect 63460 204892 63466 204904
rect 266354 204892 266360 204904
rect 266412 204892 266418 204944
rect 100754 203600 100760 203652
rect 100812 203640 100818 203652
rect 261110 203640 261116 203652
rect 100812 203612 261116 203640
rect 100812 203600 100818 203612
rect 261110 203600 261116 203612
rect 261168 203600 261174 203652
rect 155218 203532 155224 203584
rect 155276 203572 155282 203584
rect 339770 203572 339776 203584
rect 155276 203544 339776 203572
rect 155276 203532 155282 203544
rect 339770 203532 339776 203544
rect 339828 203532 339834 203584
rect 3050 202784 3056 202836
rect 3108 202824 3114 202836
rect 120074 202824 120080 202836
rect 3108 202796 120080 202824
rect 3108 202784 3114 202796
rect 120074 202784 120080 202796
rect 120132 202784 120138 202836
rect 103698 202172 103704 202224
rect 103756 202212 103762 202224
rect 216030 202212 216036 202224
rect 103756 202184 216036 202212
rect 103756 202172 103762 202184
rect 216030 202172 216036 202184
rect 216088 202172 216094 202224
rect 104894 202104 104900 202156
rect 104952 202144 104958 202156
rect 340966 202144 340972 202156
rect 104952 202116 340972 202144
rect 104952 202104 104958 202116
rect 340966 202104 340972 202116
rect 341024 202104 341030 202156
rect 59170 200744 59176 200796
rect 59228 200784 59234 200796
rect 271966 200784 271972 200796
rect 59228 200756 271972 200784
rect 59228 200744 59234 200756
rect 271966 200744 271972 200756
rect 272024 200744 272030 200796
rect 250438 199588 250444 199640
rect 250496 199628 250502 199640
rect 338390 199628 338396 199640
rect 250496 199600 338396 199628
rect 250496 199588 250502 199600
rect 338390 199588 338396 199600
rect 338448 199588 338454 199640
rect 57698 199520 57704 199572
rect 57756 199560 57762 199572
rect 258074 199560 258080 199572
rect 57756 199532 258080 199560
rect 57756 199520 57762 199532
rect 258074 199520 258080 199532
rect 258132 199520 258138 199572
rect 60550 199452 60556 199504
rect 60608 199492 60614 199504
rect 276106 199492 276112 199504
rect 60608 199464 276112 199492
rect 60608 199452 60614 199464
rect 276106 199452 276112 199464
rect 276164 199452 276170 199504
rect 87046 199384 87052 199436
rect 87104 199424 87110 199436
rect 323026 199424 323032 199436
rect 87104 199396 323032 199424
rect 87104 199384 87110 199396
rect 323026 199384 323032 199396
rect 323084 199384 323090 199436
rect 89714 198024 89720 198076
rect 89772 198064 89778 198076
rect 254210 198064 254216 198076
rect 89772 198036 254216 198064
rect 89772 198024 89778 198036
rect 254210 198024 254216 198036
rect 254268 198024 254274 198076
rect 63126 197956 63132 198008
rect 63184 197996 63190 198008
rect 262306 197996 262312 198008
rect 63184 197968 262312 197996
rect 63184 197956 63190 197968
rect 262306 197956 262312 197968
rect 262364 197956 262370 198008
rect 99466 196596 99472 196648
rect 99524 196636 99530 196648
rect 249794 196636 249800 196648
rect 99524 196608 249800 196636
rect 99524 196596 99530 196608
rect 249794 196596 249800 196608
rect 249852 196596 249858 196648
rect 86954 195304 86960 195356
rect 87012 195344 87018 195356
rect 267918 195344 267924 195356
rect 87012 195316 267924 195344
rect 87012 195304 87018 195316
rect 267918 195304 267924 195316
rect 267976 195304 267982 195356
rect 99374 195236 99380 195288
rect 99432 195276 99438 195288
rect 328638 195276 328644 195288
rect 99432 195248 328644 195276
rect 99432 195236 99438 195248
rect 328638 195236 328644 195248
rect 328696 195236 328702 195288
rect 66070 194080 66076 194132
rect 66128 194120 66134 194132
rect 251266 194120 251272 194132
rect 66128 194092 251272 194120
rect 66128 194080 66134 194092
rect 251266 194080 251272 194092
rect 251324 194080 251330 194132
rect 57514 194012 57520 194064
rect 57572 194052 57578 194064
rect 273438 194052 273444 194064
rect 57572 194024 273444 194052
rect 57572 194012 57578 194024
rect 273438 194012 273444 194024
rect 273496 194012 273502 194064
rect 65978 193944 65984 193996
rect 66036 193984 66042 193996
rect 324406 193984 324412 193996
rect 66036 193956 324412 193984
rect 66036 193944 66042 193956
rect 324406 193944 324412 193956
rect 324464 193944 324470 193996
rect 88426 193876 88432 193928
rect 88484 193916 88490 193928
rect 347866 193916 347872 193928
rect 88484 193888 347872 193916
rect 88484 193876 88490 193888
rect 347866 193876 347872 193888
rect 347924 193876 347930 193928
rect 64506 193808 64512 193860
rect 64564 193848 64570 193860
rect 347958 193848 347964 193860
rect 64564 193820 347964 193848
rect 64564 193808 64570 193820
rect 347958 193808 347964 193820
rect 348016 193808 348022 193860
rect 574738 193128 574744 193180
rect 574796 193168 574802 193180
rect 580166 193168 580172 193180
rect 574796 193140 580172 193168
rect 574796 193128 574802 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 106918 192448 106924 192500
rect 106976 192488 106982 192500
rect 259546 192488 259552 192500
rect 106976 192460 259552 192488
rect 106976 192448 106982 192460
rect 259546 192448 259552 192460
rect 259604 192448 259610 192500
rect 92566 191360 92572 191412
rect 92624 191400 92630 191412
rect 249886 191400 249892 191412
rect 92624 191372 249892 191400
rect 92624 191360 92630 191372
rect 249886 191360 249892 191372
rect 249944 191360 249950 191412
rect 84194 191292 84200 191344
rect 84252 191332 84258 191344
rect 321738 191332 321744 191344
rect 84252 191304 321744 191332
rect 84252 191292 84258 191304
rect 321738 191292 321744 191304
rect 321796 191292 321802 191344
rect 107654 191224 107660 191276
rect 107712 191264 107718 191276
rect 347774 191264 347780 191276
rect 107712 191236 347780 191264
rect 107712 191224 107718 191236
rect 347774 191224 347780 191236
rect 347832 191224 347838 191276
rect 95326 191156 95332 191208
rect 95384 191196 95390 191208
rect 336826 191196 336832 191208
rect 95384 191168 336832 191196
rect 95384 191156 95390 191168
rect 336826 191156 336832 191168
rect 336884 191156 336890 191208
rect 102134 191088 102140 191140
rect 102192 191128 102198 191140
rect 343910 191128 343916 191140
rect 102192 191100 343916 191128
rect 102192 191088 102198 191100
rect 343910 191088 343916 191100
rect 343968 191088 343974 191140
rect 169018 189796 169024 189848
rect 169076 189836 169082 189848
rect 269206 189836 269212 189848
rect 169076 189808 269212 189836
rect 169076 189796 169082 189808
rect 269206 189796 269212 189808
rect 269264 189796 269270 189848
rect 73154 189728 73160 189780
rect 73212 189768 73218 189780
rect 325878 189768 325884 189780
rect 73212 189740 325884 189768
rect 73212 189728 73218 189740
rect 325878 189728 325884 189740
rect 325936 189728 325942 189780
rect 106182 189048 106188 189100
rect 106240 189088 106246 189100
rect 173158 189088 173164 189100
rect 106240 189060 173164 189088
rect 106240 189048 106246 189060
rect 173158 189048 173164 189060
rect 173216 189048 173222 189100
rect 160738 188572 160744 188624
rect 160796 188612 160802 188624
rect 274726 188612 274732 188624
rect 160796 188584 274732 188612
rect 160796 188572 160802 188584
rect 274726 188572 274732 188584
rect 274784 188572 274790 188624
rect 214650 188504 214656 188556
rect 214708 188544 214714 188556
rect 334158 188544 334164 188556
rect 214708 188516 334164 188544
rect 214708 188504 214714 188516
rect 334158 188504 334164 188516
rect 334216 188504 334222 188556
rect 55030 188436 55036 188488
rect 55088 188476 55094 188488
rect 259638 188476 259644 188488
rect 55088 188448 259644 188476
rect 55088 188436 55094 188448
rect 259638 188436 259644 188448
rect 259696 188436 259702 188488
rect 64782 188368 64788 188420
rect 64840 188408 64846 188420
rect 270586 188408 270592 188420
rect 64840 188380 270592 188408
rect 64840 188368 64846 188380
rect 270586 188368 270592 188380
rect 270644 188368 270650 188420
rect 70394 188300 70400 188352
rect 70452 188340 70458 188352
rect 345198 188340 345204 188352
rect 70452 188312 345204 188340
rect 70452 188300 70458 188312
rect 345198 188300 345204 188312
rect 345256 188300 345262 188352
rect 107562 187756 107568 187808
rect 107620 187796 107626 187808
rect 171778 187796 171784 187808
rect 107620 187768 171784 187796
rect 107620 187756 107626 187768
rect 171778 187756 171784 187768
rect 171836 187756 171842 187808
rect 133782 187688 133788 187740
rect 133840 187728 133846 187740
rect 214558 187728 214564 187740
rect 133840 187700 214564 187728
rect 133840 187688 133846 187700
rect 214558 187688 214564 187700
rect 214616 187688 214622 187740
rect 206278 187008 206284 187060
rect 206336 187048 206342 187060
rect 274634 187048 274640 187060
rect 206336 187020 274640 187048
rect 206336 187008 206342 187020
rect 274634 187008 274640 187020
rect 274692 187008 274698 187060
rect 17218 186940 17224 186992
rect 17276 186980 17282 186992
rect 110414 186980 110420 186992
rect 17276 186952 110420 186980
rect 17276 186940 17282 186952
rect 110414 186940 110420 186952
rect 110472 186940 110478 186992
rect 152458 186940 152464 186992
rect 152516 186980 152522 186992
rect 331306 186980 331312 186992
rect 152516 186952 331312 186980
rect 152516 186940 152522 186952
rect 331306 186940 331312 186952
rect 331364 186940 331370 186992
rect 132402 186464 132408 186516
rect 132460 186504 132466 186516
rect 170582 186504 170588 186516
rect 132460 186476 170588 186504
rect 132460 186464 132466 186476
rect 170582 186464 170588 186476
rect 170640 186464 170646 186516
rect 100662 186396 100668 186448
rect 100720 186436 100726 186448
rect 169018 186436 169024 186448
rect 100720 186408 169024 186436
rect 100720 186396 100726 186408
rect 169018 186396 169024 186408
rect 169076 186396 169082 186448
rect 118602 186328 118608 186380
rect 118660 186368 118666 186380
rect 214650 186368 214656 186380
rect 118660 186340 214656 186368
rect 118660 186328 118666 186340
rect 214650 186328 214656 186340
rect 214708 186328 214714 186380
rect 118694 185852 118700 185904
rect 118752 185892 118758 185904
rect 346578 185892 346584 185904
rect 118752 185864 346584 185892
rect 118752 185852 118758 185864
rect 346578 185852 346584 185864
rect 346636 185852 346642 185904
rect 80054 185784 80060 185836
rect 80112 185824 80118 185836
rect 327350 185824 327356 185836
rect 80112 185796 327356 185824
rect 80112 185784 80118 185796
rect 327350 185784 327356 185796
rect 327408 185784 327414 185836
rect 65886 185716 65892 185768
rect 65944 185756 65950 185768
rect 324498 185756 324504 185768
rect 65944 185728 324504 185756
rect 65944 185716 65950 185728
rect 324498 185716 324504 185728
rect 324556 185716 324562 185768
rect 67542 185648 67548 185700
rect 67600 185688 67606 185700
rect 334250 185688 334256 185700
rect 67600 185660 334256 185688
rect 67600 185648 67606 185660
rect 334250 185648 334256 185660
rect 334308 185648 334314 185700
rect 58986 185580 58992 185632
rect 59044 185620 59050 185632
rect 331398 185620 331404 185632
rect 59044 185592 331404 185620
rect 59044 185580 59050 185592
rect 331398 185580 331404 185592
rect 331456 185580 331462 185632
rect 121362 184900 121368 184952
rect 121420 184940 121426 184952
rect 170490 184940 170496 184952
rect 121420 184912 170496 184940
rect 121420 184900 121426 184912
rect 170490 184900 170496 184912
rect 170548 184900 170554 184952
rect 180058 184288 180064 184340
rect 180116 184328 180122 184340
rect 262398 184328 262404 184340
rect 180116 184300 262404 184328
rect 180116 184288 180122 184300
rect 262398 184288 262404 184300
rect 262456 184288 262462 184340
rect 289078 184288 289084 184340
rect 289136 184328 289142 184340
rect 338206 184328 338212 184340
rect 289136 184300 338212 184328
rect 289136 184288 289142 184300
rect 338206 184288 338212 184300
rect 338264 184288 338270 184340
rect 57790 184220 57796 184272
rect 57848 184260 57854 184272
rect 308490 184260 308496 184272
rect 57848 184232 308496 184260
rect 57848 184220 57854 184232
rect 308490 184220 308496 184232
rect 308548 184220 308554 184272
rect 69014 184152 69020 184204
rect 69072 184192 69078 184204
rect 323210 184192 323216 184204
rect 69072 184164 323216 184192
rect 69072 184152 69078 184164
rect 323210 184152 323216 184164
rect 323268 184152 323274 184204
rect 114462 183540 114468 183592
rect 114520 183580 114526 183592
rect 169294 183580 169300 183592
rect 114520 183552 169300 183580
rect 114520 183540 114526 183552
rect 169294 183540 169300 183552
rect 169352 183540 169358 183592
rect 244918 183132 244924 183184
rect 244976 183172 244982 183184
rect 256786 183172 256792 183184
rect 244976 183144 256792 183172
rect 244976 183132 244982 183144
rect 256786 183132 256792 183144
rect 256844 183132 256850 183184
rect 238110 183064 238116 183116
rect 238168 183104 238174 183116
rect 256970 183104 256976 183116
rect 238168 183076 256976 183104
rect 238168 183064 238174 183076
rect 256970 183064 256976 183076
rect 257028 183064 257034 183116
rect 213178 182996 213184 183048
rect 213236 183036 213242 183048
rect 265066 183036 265072 183048
rect 213236 183008 265072 183036
rect 213236 182996 213242 183008
rect 265066 182996 265072 183008
rect 265124 182996 265130 183048
rect 186958 182928 186964 182980
rect 187016 182968 187022 182980
rect 262490 182968 262496 182980
rect 187016 182940 262496 182968
rect 187016 182928 187022 182940
rect 262490 182928 262496 182940
rect 262548 182928 262554 182980
rect 276658 182928 276664 182980
rect 276716 182968 276722 182980
rect 336918 182968 336924 182980
rect 276716 182940 336924 182968
rect 276716 182928 276722 182940
rect 336918 182928 336924 182940
rect 336976 182928 336982 182980
rect 93854 182860 93860 182912
rect 93912 182900 93918 182912
rect 338482 182900 338488 182912
rect 93912 182872 338488 182900
rect 93912 182860 93918 182872
rect 338482 182860 338488 182872
rect 338540 182860 338546 182912
rect 56502 182792 56508 182844
rect 56560 182832 56566 182844
rect 345290 182832 345296 182844
rect 56560 182804 345296 182832
rect 56560 182792 56566 182804
rect 345290 182792 345296 182804
rect 345348 182792 345354 182844
rect 116946 182316 116952 182368
rect 117004 182356 117010 182368
rect 167730 182356 167736 182368
rect 117004 182328 167736 182356
rect 117004 182316 117010 182328
rect 167730 182316 167736 182328
rect 167788 182316 167794 182368
rect 97534 182248 97540 182300
rect 97592 182288 97598 182300
rect 169202 182288 169208 182300
rect 97592 182260 169208 182288
rect 97592 182248 97598 182260
rect 169202 182248 169208 182260
rect 169260 182248 169266 182300
rect 129458 182180 129464 182232
rect 129516 182220 129522 182232
rect 213270 182220 213276 182232
rect 129516 182192 213276 182220
rect 129516 182180 129522 182192
rect 213270 182180 213276 182192
rect 213328 182180 213334 182232
rect 316678 181636 316684 181688
rect 316736 181676 316742 181688
rect 342530 181676 342536 181688
rect 316736 181648 342536 181676
rect 316736 181636 316742 181648
rect 342530 181636 342536 181648
rect 342588 181636 342594 181688
rect 202138 181568 202144 181620
rect 202196 181608 202202 181620
rect 246942 181608 246948 181620
rect 202196 181580 246948 181608
rect 202196 181568 202202 181580
rect 246942 181568 246948 181580
rect 247000 181568 247006 181620
rect 300118 181568 300124 181620
rect 300176 181608 300182 181620
rect 332686 181608 332692 181620
rect 300176 181580 332692 181608
rect 300176 181568 300182 181580
rect 332686 181568 332692 181580
rect 332744 181568 332750 181620
rect 170398 181500 170404 181552
rect 170456 181540 170462 181552
rect 316310 181540 316316 181552
rect 170456 181512 316316 181540
rect 170456 181500 170462 181512
rect 316310 181500 316316 181512
rect 316368 181500 316374 181552
rect 318058 181500 318064 181552
rect 318116 181540 318122 181552
rect 341150 181540 341156 181552
rect 318116 181512 341156 181540
rect 318116 181500 318122 181512
rect 341150 181500 341156 181512
rect 341208 181500 341214 181552
rect 74718 181432 74724 181484
rect 74776 181472 74782 181484
rect 252830 181472 252836 181484
rect 74776 181444 252836 181472
rect 74776 181432 74782 181444
rect 252830 181432 252836 181444
rect 252888 181432 252894 181484
rect 307018 181432 307024 181484
rect 307076 181472 307082 181484
rect 339678 181472 339684 181484
rect 307076 181444 339684 181472
rect 307076 181432 307082 181444
rect 339678 181432 339684 181444
rect 339736 181432 339742 181484
rect 112990 180820 112996 180872
rect 113048 180860 113054 180872
rect 166350 180860 166356 180872
rect 113048 180832 166356 180860
rect 113048 180820 113054 180832
rect 166350 180820 166356 180832
rect 166408 180820 166414 180872
rect 238018 180412 238024 180464
rect 238076 180452 238082 180464
rect 261018 180452 261024 180464
rect 238076 180424 261024 180452
rect 238076 180412 238082 180424
rect 261018 180412 261024 180424
rect 261076 180412 261082 180464
rect 228358 180344 228364 180396
rect 228416 180384 228422 180396
rect 259454 180384 259460 180396
rect 228416 180356 259460 180384
rect 228416 180344 228422 180356
rect 259454 180344 259460 180356
rect 259512 180344 259518 180396
rect 222838 180276 222844 180328
rect 222896 180316 222902 180328
rect 258166 180316 258172 180328
rect 222896 180288 258172 180316
rect 222896 180276 222902 180288
rect 258166 180276 258172 180288
rect 258224 180276 258230 180328
rect 191190 180208 191196 180260
rect 191248 180248 191254 180260
rect 255590 180248 255596 180260
rect 191248 180220 255596 180248
rect 191248 180208 191254 180220
rect 255590 180208 255596 180220
rect 255648 180208 255654 180260
rect 72418 180140 72424 180192
rect 72476 180180 72482 180192
rect 332778 180180 332784 180192
rect 72476 180152 332784 180180
rect 72476 180140 72482 180152
rect 332778 180140 332784 180152
rect 332836 180140 332842 180192
rect 67450 180072 67456 180124
rect 67508 180112 67514 180124
rect 335538 180112 335544 180124
rect 67508 180084 335544 180112
rect 67508 180072 67514 180084
rect 335538 180072 335544 180084
rect 335596 180072 335602 180124
rect 123754 179460 123760 179512
rect 123812 179500 123818 179512
rect 167822 179500 167828 179512
rect 123812 179472 167828 179500
rect 123812 179460 123818 179472
rect 167822 179460 167828 179472
rect 167880 179460 167886 179512
rect 128078 179392 128084 179444
rect 128136 179432 128142 179444
rect 211798 179432 211804 179444
rect 128136 179404 211804 179432
rect 128136 179392 128142 179404
rect 211798 179392 211804 179404
rect 211856 179392 211862 179444
rect 287698 179324 287704 179376
rect 287756 179364 287762 179376
rect 338298 179364 338304 179376
rect 287756 179336 338304 179364
rect 287756 179324 287762 179336
rect 338298 179324 338304 179336
rect 338356 179324 338362 179376
rect 231118 178916 231124 178968
rect 231176 178956 231182 178968
rect 249058 178956 249064 178968
rect 231176 178928 249064 178956
rect 231176 178916 231182 178928
rect 249058 178916 249064 178928
rect 249116 178916 249122 178968
rect 209038 178848 209044 178900
rect 209096 178888 209102 178900
rect 249242 178888 249248 178900
rect 209096 178860 249248 178888
rect 209096 178848 209102 178860
rect 249242 178848 249248 178860
rect 249300 178848 249306 178900
rect 215938 178780 215944 178832
rect 215996 178820 216002 178832
rect 258258 178820 258264 178832
rect 215996 178792 258264 178820
rect 215996 178780 216002 178792
rect 258258 178780 258264 178792
rect 258316 178780 258322 178832
rect 204898 178712 204904 178764
rect 204956 178752 204962 178764
rect 260834 178752 260840 178764
rect 204956 178724 260840 178752
rect 204956 178712 204962 178724
rect 260834 178712 260840 178724
rect 260892 178712 260898 178764
rect 162118 178644 162124 178696
rect 162176 178684 162182 178696
rect 331490 178684 331496 178696
rect 162176 178656 331496 178684
rect 162176 178644 162182 178656
rect 331490 178644 331496 178656
rect 331548 178644 331554 178696
rect 148226 178304 148232 178356
rect 148284 178344 148290 178356
rect 169110 178344 169116 178356
rect 148284 178316 169116 178344
rect 148284 178304 148290 178316
rect 169110 178304 169116 178316
rect 169168 178304 169174 178356
rect 134794 178236 134800 178288
rect 134852 178276 134858 178288
rect 165338 178276 165344 178288
rect 134852 178248 165344 178276
rect 134852 178236 134858 178248
rect 165338 178236 165344 178248
rect 165396 178236 165402 178288
rect 126054 178168 126060 178220
rect 126112 178208 126118 178220
rect 167914 178208 167920 178220
rect 126112 178180 167920 178208
rect 126112 178168 126118 178180
rect 167914 178168 167920 178180
rect 167972 178168 167978 178220
rect 115842 178100 115848 178152
rect 115900 178140 115906 178152
rect 166442 178140 166448 178152
rect 115900 178112 166448 178140
rect 115900 178100 115906 178112
rect 166442 178100 166448 178112
rect 166500 178100 166506 178152
rect 109954 178032 109960 178084
rect 110012 178072 110018 178084
rect 170398 178072 170404 178084
rect 110012 178044 170404 178072
rect 110012 178032 110018 178044
rect 170398 178032 170404 178044
rect 170456 178032 170462 178084
rect 242158 177964 242164 178016
rect 242216 178004 242222 178016
rect 249150 178004 249156 178016
rect 242216 177976 249156 178004
rect 242216 177964 242222 177976
rect 249150 177964 249156 177976
rect 249208 177964 249214 178016
rect 312538 177488 312544 177540
rect 312596 177528 312602 177540
rect 332594 177528 332600 177540
rect 312596 177500 332600 177528
rect 312596 177488 312602 177500
rect 332594 177488 332600 177500
rect 332652 177488 332658 177540
rect 246298 177420 246304 177472
rect 246356 177460 246362 177472
rect 263778 177460 263784 177472
rect 246356 177432 263784 177460
rect 246356 177420 246362 177432
rect 263778 177420 263784 177432
rect 263836 177420 263842 177472
rect 315298 177420 315304 177472
rect 315356 177460 315362 177472
rect 335630 177460 335636 177472
rect 315356 177432 335636 177460
rect 315356 177420 315362 177432
rect 335630 177420 335636 177432
rect 335688 177420 335694 177472
rect 233970 177352 233976 177404
rect 234028 177392 234034 177404
rect 258350 177392 258356 177404
rect 234028 177364 258356 177392
rect 234028 177352 234034 177364
rect 258350 177352 258356 177364
rect 258408 177352 258414 177404
rect 304258 177352 304264 177404
rect 304316 177392 304322 177404
rect 333974 177392 333980 177404
rect 304316 177364 333980 177392
rect 304316 177352 304322 177364
rect 333974 177352 333980 177364
rect 334032 177352 334038 177404
rect 4798 177284 4804 177336
rect 4856 177324 4862 177336
rect 82814 177324 82820 177336
rect 4856 177296 82820 177324
rect 4856 177284 4862 177296
rect 82814 177284 82820 177296
rect 82872 177284 82878 177336
rect 195238 177284 195244 177336
rect 195296 177324 195302 177336
rect 251358 177324 251364 177336
rect 195296 177296 251364 177324
rect 195296 177284 195302 177296
rect 251358 177284 251364 177296
rect 251416 177284 251422 177336
rect 284938 177284 284944 177336
rect 284996 177324 285002 177336
rect 337010 177324 337016 177336
rect 284996 177296 337016 177324
rect 284996 177284 285002 177296
rect 337010 177284 337016 177296
rect 337068 177284 337074 177336
rect 130746 177012 130752 177064
rect 130804 177052 130810 177064
rect 165522 177052 165528 177064
rect 130804 177024 165528 177052
rect 130804 177012 130810 177024
rect 165522 177012 165528 177024
rect 165580 177012 165586 177064
rect 104618 176944 104624 176996
rect 104676 176984 104682 176996
rect 165430 176984 165436 176996
rect 104676 176956 165436 176984
rect 104676 176944 104682 176956
rect 165430 176944 165436 176956
rect 165488 176944 165494 176996
rect 103330 176876 103336 176928
rect 103388 176916 103394 176928
rect 167638 176916 167644 176928
rect 103388 176888 167644 176916
rect 103388 176876 103394 176888
rect 167638 176876 167644 176888
rect 167696 176876 167702 176928
rect 136082 176808 136088 176860
rect 136140 176848 136146 176860
rect 213914 176848 213920 176860
rect 136140 176820 213920 176848
rect 136140 176808 136146 176820
rect 213914 176808 213920 176820
rect 213972 176808 213978 176860
rect 124490 176740 124496 176792
rect 124548 176780 124554 176792
rect 211890 176780 211896 176792
rect 124548 176752 211896 176780
rect 124548 176740 124554 176752
rect 211890 176740 211896 176752
rect 211948 176740 211954 176792
rect 108114 176672 108120 176724
rect 108172 176712 108178 176724
rect 195330 176712 195336 176724
rect 108172 176684 195336 176712
rect 108172 176672 108178 176684
rect 195330 176672 195336 176684
rect 195388 176672 195394 176724
rect 305638 176604 305644 176656
rect 305696 176644 305702 176656
rect 321462 176644 321468 176656
rect 305696 176616 321468 176644
rect 305696 176604 305702 176616
rect 321462 176604 321468 176616
rect 321520 176604 321526 176656
rect 158898 176264 158904 176316
rect 158956 176304 158962 176316
rect 166258 176304 166264 176316
rect 158956 176276 166264 176304
rect 158956 176264 158962 176276
rect 166258 176264 166264 176276
rect 166316 176264 166322 176316
rect 121914 176196 121920 176248
rect 121972 176236 121978 176248
rect 166534 176236 166540 176248
rect 121972 176208 166540 176236
rect 121972 176196 121978 176208
rect 166534 176196 166540 176208
rect 166592 176196 166598 176248
rect 113174 176128 113180 176180
rect 113232 176168 113238 176180
rect 170674 176168 170680 176180
rect 113232 176140 170680 176168
rect 113232 176128 113238 176140
rect 170674 176128 170680 176140
rect 170732 176128 170738 176180
rect 128170 176060 128176 176112
rect 128228 176100 128234 176112
rect 212258 176100 212264 176112
rect 128228 176072 212264 176100
rect 128228 176060 128234 176072
rect 212258 176060 212264 176072
rect 212316 176060 212322 176112
rect 119430 175992 119436 176044
rect 119488 176032 119494 176044
rect 214742 176032 214748 176044
rect 119488 176004 214748 176032
rect 119488 175992 119494 176004
rect 214742 175992 214748 176004
rect 214800 175992 214806 176044
rect 240778 175992 240784 176044
rect 240836 176032 240842 176044
rect 256694 176032 256700 176044
rect 240836 176004 256700 176032
rect 240836 175992 240842 176004
rect 256694 175992 256700 176004
rect 256752 175992 256758 176044
rect 338390 175992 338396 176044
rect 338448 175992 338454 176044
rect 100754 175924 100760 175976
rect 100812 175964 100818 175976
rect 209038 175964 209044 175976
rect 100812 175936 209044 175964
rect 100812 175924 100818 175936
rect 209038 175924 209044 175936
rect 209096 175924 209102 175976
rect 233878 175924 233884 175976
rect 233936 175964 233942 175976
rect 249978 175964 249984 175976
rect 233936 175936 249984 175964
rect 233936 175924 233942 175936
rect 249978 175924 249984 175936
rect 250036 175924 250042 175976
rect 313918 175924 313924 175976
rect 313976 175964 313982 175976
rect 321462 175964 321468 175976
rect 313976 175936 321468 175964
rect 313976 175924 313982 175936
rect 321462 175924 321468 175936
rect 321520 175924 321526 175976
rect 338408 175840 338436 175992
rect 338390 175788 338396 175840
rect 338448 175788 338454 175840
rect 165338 175176 165344 175228
rect 165396 175216 165402 175228
rect 213914 175216 213920 175228
rect 165396 175188 213920 175216
rect 165396 175176 165402 175188
rect 213914 175176 213920 175188
rect 213972 175176 213978 175228
rect 165522 174496 165528 174548
rect 165580 174536 165586 174548
rect 214006 174536 214012 174548
rect 165580 174508 214012 174536
rect 165580 174496 165586 174508
rect 214006 174496 214012 174508
rect 214064 174496 214070 174548
rect 287790 174020 287796 174072
rect 287848 174060 287854 174072
rect 307570 174060 307576 174072
rect 287848 174032 307576 174060
rect 287848 174020 287854 174032
rect 307570 174020 307576 174032
rect 307628 174020 307634 174072
rect 268378 173952 268384 174004
rect 268436 173992 268442 174004
rect 307662 173992 307668 174004
rect 268436 173964 307668 173992
rect 268436 173952 268442 173964
rect 307662 173952 307668 173964
rect 307720 173952 307726 174004
rect 264238 173884 264244 173936
rect 264296 173924 264302 173936
rect 306558 173924 306564 173936
rect 264296 173896 306564 173924
rect 264296 173884 264302 173896
rect 306558 173884 306564 173896
rect 306616 173884 306622 173936
rect 170582 173816 170588 173868
rect 170640 173856 170646 173868
rect 213914 173856 213920 173868
rect 170640 173828 213920 173856
rect 170640 173816 170646 173828
rect 213914 173816 213920 173828
rect 213972 173816 213978 173868
rect 165430 173136 165436 173188
rect 165488 173176 165494 173188
rect 214650 173176 214656 173188
rect 165488 173148 214656 173176
rect 165488 173136 165494 173148
rect 214650 173136 214656 173148
rect 214708 173136 214714 173188
rect 284938 172660 284944 172712
rect 284996 172700 285002 172712
rect 307478 172700 307484 172712
rect 284996 172672 307484 172700
rect 284996 172660 285002 172672
rect 307478 172660 307484 172672
rect 307536 172660 307542 172712
rect 276658 172592 276664 172644
rect 276716 172632 276722 172644
rect 307570 172632 307576 172644
rect 276716 172604 307576 172632
rect 276716 172592 276722 172604
rect 307570 172592 307576 172604
rect 307628 172592 307634 172644
rect 252462 172524 252468 172576
rect 252520 172564 252526 172576
rect 259638 172564 259644 172576
rect 252520 172536 259644 172564
rect 252520 172524 252526 172536
rect 259638 172524 259644 172536
rect 259696 172524 259702 172576
rect 267182 172524 267188 172576
rect 267240 172564 267246 172576
rect 307662 172564 307668 172576
rect 267240 172536 307668 172564
rect 267240 172524 267246 172536
rect 307662 172524 307668 172536
rect 307720 172524 307726 172576
rect 212258 172456 212264 172508
rect 212316 172496 212322 172508
rect 213914 172496 213920 172508
rect 212316 172468 213920 172496
rect 212316 172456 212322 172468
rect 213914 172456 213920 172468
rect 213972 172456 213978 172508
rect 324314 172456 324320 172508
rect 324372 172496 324378 172508
rect 336826 172496 336832 172508
rect 324372 172468 336832 172496
rect 324372 172456 324378 172468
rect 336826 172456 336832 172468
rect 336884 172456 336890 172508
rect 252462 172320 252468 172372
rect 252520 172360 252526 172372
rect 263594 172360 263600 172372
rect 252520 172332 263600 172360
rect 252520 172320 252526 172332
rect 263594 172320 263600 172332
rect 263652 172320 263658 172372
rect 252370 171368 252376 171420
rect 252428 171408 252434 171420
rect 259454 171408 259460 171420
rect 252428 171380 259460 171408
rect 252428 171368 252434 171380
rect 259454 171368 259460 171380
rect 259512 171368 259518 171420
rect 289170 171232 289176 171284
rect 289228 171272 289234 171284
rect 306558 171272 306564 171284
rect 289228 171244 306564 171272
rect 289228 171232 289234 171244
rect 306558 171232 306564 171244
rect 306616 171232 306622 171284
rect 265802 171164 265808 171216
rect 265860 171204 265866 171216
rect 307570 171204 307576 171216
rect 265860 171176 307576 171204
rect 265860 171164 265866 171176
rect 307570 171164 307576 171176
rect 307628 171164 307634 171216
rect 168006 171096 168012 171148
rect 168064 171136 168070 171148
rect 214466 171136 214472 171148
rect 168064 171108 214472 171136
rect 168064 171096 168070 171108
rect 214466 171096 214472 171108
rect 214524 171096 214530 171148
rect 260282 171096 260288 171148
rect 260340 171136 260346 171148
rect 307662 171136 307668 171148
rect 260340 171108 307668 171136
rect 260340 171096 260346 171108
rect 307662 171096 307668 171108
rect 307720 171096 307726 171148
rect 167914 171028 167920 171080
rect 167972 171068 167978 171080
rect 213914 171068 213920 171080
rect 167972 171040 213920 171068
rect 167972 171028 167978 171040
rect 213914 171028 213920 171040
rect 213972 171028 213978 171080
rect 324314 171028 324320 171080
rect 324372 171068 324378 171080
rect 338114 171068 338120 171080
rect 324372 171040 338120 171068
rect 324372 171028 324378 171040
rect 338114 171028 338120 171040
rect 338172 171028 338178 171080
rect 211798 170960 211804 171012
rect 211856 171000 211862 171012
rect 214466 171000 214472 171012
rect 211856 170972 214472 171000
rect 211856 170960 211862 170972
rect 214466 170960 214472 170972
rect 214524 170960 214530 171012
rect 252462 170756 252468 170808
rect 252520 170796 252526 170808
rect 256694 170796 256700 170808
rect 252520 170768 256700 170796
rect 252520 170756 252526 170768
rect 256694 170756 256700 170768
rect 256752 170756 256758 170808
rect 286410 169872 286416 169924
rect 286468 169912 286474 169924
rect 306558 169912 306564 169924
rect 286468 169884 306564 169912
rect 286468 169872 286474 169884
rect 306558 169872 306564 169884
rect 306616 169872 306622 169924
rect 252462 169804 252468 169856
rect 252520 169844 252526 169856
rect 258074 169844 258080 169856
rect 252520 169816 258080 169844
rect 252520 169804 252526 169816
rect 258074 169804 258080 169816
rect 258132 169804 258138 169856
rect 265710 169804 265716 169856
rect 265768 169844 265774 169856
rect 307570 169844 307576 169856
rect 265768 169816 307576 169844
rect 265768 169804 265774 169816
rect 307570 169804 307576 169816
rect 307628 169804 307634 169856
rect 258994 169736 259000 169788
rect 259052 169776 259058 169788
rect 307662 169776 307668 169788
rect 259052 169748 307668 169776
rect 259052 169736 259058 169748
rect 307662 169736 307668 169748
rect 307720 169736 307726 169788
rect 167822 169668 167828 169720
rect 167880 169708 167886 169720
rect 213914 169708 213920 169720
rect 167880 169680 213920 169708
rect 167880 169668 167886 169680
rect 213914 169668 213920 169680
rect 213972 169668 213978 169720
rect 252370 169668 252376 169720
rect 252428 169708 252434 169720
rect 260926 169708 260932 169720
rect 252428 169680 260932 169708
rect 252428 169668 252434 169680
rect 260926 169668 260932 169680
rect 260984 169668 260990 169720
rect 211890 169600 211896 169652
rect 211948 169640 211954 169652
rect 214006 169640 214012 169652
rect 211948 169612 214012 169640
rect 211948 169600 211954 169612
rect 214006 169600 214012 169612
rect 214064 169600 214070 169652
rect 252278 169600 252284 169652
rect 252336 169640 252342 169652
rect 260834 169640 260840 169652
rect 252336 169612 260840 169640
rect 252336 169600 252342 169612
rect 260834 169600 260840 169612
rect 260892 169600 260898 169652
rect 252462 168920 252468 168972
rect 252520 168960 252526 168972
rect 259546 168960 259552 168972
rect 252520 168932 259552 168960
rect 252520 168920 252526 168932
rect 259546 168920 259552 168932
rect 259604 168920 259610 168972
rect 291838 168512 291844 168564
rect 291896 168552 291902 168564
rect 307662 168552 307668 168564
rect 291896 168524 307668 168552
rect 291896 168512 291902 168524
rect 307662 168512 307668 168524
rect 307720 168512 307726 168564
rect 269850 168444 269856 168496
rect 269908 168484 269914 168496
rect 307478 168484 307484 168496
rect 269908 168456 307484 168484
rect 269908 168444 269914 168456
rect 307478 168444 307484 168456
rect 307536 168444 307542 168496
rect 261570 168376 261576 168428
rect 261628 168416 261634 168428
rect 307570 168416 307576 168428
rect 261628 168388 307576 168416
rect 261628 168376 261634 168388
rect 307570 168376 307576 168388
rect 307628 168376 307634 168428
rect 166534 168308 166540 168360
rect 166592 168348 166598 168360
rect 213914 168348 213920 168360
rect 166592 168320 213920 168348
rect 166592 168308 166598 168320
rect 213914 168308 213920 168320
rect 213972 168308 213978 168360
rect 252370 168308 252376 168360
rect 252428 168348 252434 168360
rect 261018 168348 261024 168360
rect 252428 168320 261024 168348
rect 252428 168308 252434 168320
rect 261018 168308 261024 168320
rect 261076 168308 261082 168360
rect 324314 168308 324320 168360
rect 324372 168348 324378 168360
rect 332778 168348 332784 168360
rect 324372 168320 332784 168348
rect 324372 168308 324378 168320
rect 332778 168308 332784 168320
rect 332836 168308 332842 168360
rect 170490 168240 170496 168292
rect 170548 168280 170554 168292
rect 214006 168280 214012 168292
rect 170548 168252 214012 168280
rect 170548 168240 170554 168252
rect 214006 168240 214012 168252
rect 214064 168240 214070 168292
rect 252278 168240 252284 168292
rect 252336 168280 252342 168292
rect 255406 168280 255412 168292
rect 252336 168252 255412 168280
rect 252336 168240 252342 168252
rect 255406 168240 255412 168252
rect 255464 168240 255470 168292
rect 324406 168240 324412 168292
rect 324464 168280 324470 168292
rect 332594 168280 332600 168292
rect 324464 168252 332600 168280
rect 324464 168240 324470 168252
rect 332594 168240 332600 168252
rect 332652 168240 332658 168292
rect 252462 167832 252468 167884
rect 252520 167872 252526 167884
rect 258258 167872 258264 167884
rect 252520 167844 258264 167872
rect 252520 167832 252526 167844
rect 258258 167832 258264 167844
rect 258316 167832 258322 167884
rect 282270 167152 282276 167204
rect 282328 167192 282334 167204
rect 307662 167192 307668 167204
rect 282328 167164 307668 167192
rect 282328 167152 282334 167164
rect 307662 167152 307668 167164
rect 307720 167152 307726 167204
rect 271322 167084 271328 167136
rect 271380 167124 271386 167136
rect 307570 167124 307576 167136
rect 271380 167096 307576 167124
rect 271380 167084 271386 167096
rect 307570 167084 307576 167096
rect 307628 167084 307634 167136
rect 261662 167016 261668 167068
rect 261720 167056 261726 167068
rect 307478 167056 307484 167068
rect 261720 167028 307484 167056
rect 261720 167016 261726 167028
rect 307478 167016 307484 167028
rect 307536 167016 307542 167068
rect 167730 166948 167736 167000
rect 167788 166988 167794 167000
rect 213914 166988 213920 167000
rect 167788 166960 213920 166988
rect 167788 166948 167794 166960
rect 213914 166948 213920 166960
rect 213972 166948 213978 167000
rect 324314 166948 324320 167000
rect 324372 166988 324378 167000
rect 335630 166988 335636 167000
rect 324372 166960 335636 166988
rect 324372 166948 324378 166960
rect 335630 166948 335636 166960
rect 335688 166948 335694 167000
rect 252462 166200 252468 166252
rect 252520 166240 252526 166252
rect 258166 166240 258172 166252
rect 252520 166212 258172 166240
rect 252520 166200 252526 166212
rect 258166 166200 258172 166212
rect 258224 166200 258230 166252
rect 252370 165724 252376 165776
rect 252428 165764 252434 165776
rect 258350 165764 258356 165776
rect 252428 165736 258356 165764
rect 252428 165724 252434 165736
rect 258350 165724 258356 165736
rect 258408 165724 258414 165776
rect 280798 165724 280804 165776
rect 280856 165764 280862 165776
rect 307662 165764 307668 165776
rect 280856 165736 307668 165764
rect 280856 165724 280862 165736
rect 307662 165724 307668 165736
rect 307720 165724 307726 165776
rect 272610 165656 272616 165708
rect 272668 165696 272674 165708
rect 307294 165696 307300 165708
rect 272668 165668 307300 165696
rect 272668 165656 272674 165668
rect 307294 165656 307300 165668
rect 307352 165656 307358 165708
rect 258902 165588 258908 165640
rect 258960 165628 258966 165640
rect 307570 165628 307576 165640
rect 258960 165600 307576 165628
rect 258960 165588 258966 165600
rect 307570 165588 307576 165600
rect 307628 165588 307634 165640
rect 166442 165520 166448 165572
rect 166500 165560 166506 165572
rect 213914 165560 213920 165572
rect 166500 165532 213920 165560
rect 166500 165520 166506 165532
rect 213914 165520 213920 165532
rect 213972 165520 213978 165572
rect 252370 165520 252376 165572
rect 252428 165560 252434 165572
rect 264974 165560 264980 165572
rect 252428 165532 264980 165560
rect 252428 165520 252434 165532
rect 264974 165520 264980 165532
rect 265032 165520 265038 165572
rect 324314 165520 324320 165572
rect 324372 165560 324378 165572
rect 343910 165560 343916 165572
rect 324372 165532 343916 165560
rect 324372 165520 324378 165532
rect 343910 165520 343916 165532
rect 343968 165520 343974 165572
rect 169294 165452 169300 165504
rect 169352 165492 169358 165504
rect 214006 165492 214012 165504
rect 169352 165464 214012 165492
rect 169352 165452 169358 165464
rect 214006 165452 214012 165464
rect 214064 165452 214070 165504
rect 252462 165452 252468 165504
rect 252520 165492 252526 165504
rect 262490 165492 262496 165504
rect 252520 165464 262496 165492
rect 252520 165452 252526 165464
rect 262490 165452 262496 165464
rect 262548 165452 262554 165504
rect 300394 164364 300400 164416
rect 300452 164404 300458 164416
rect 307570 164404 307576 164416
rect 300452 164376 307576 164404
rect 300452 164364 300458 164376
rect 307570 164364 307576 164376
rect 307628 164364 307634 164416
rect 274082 164296 274088 164348
rect 274140 164336 274146 164348
rect 307662 164336 307668 164348
rect 274140 164308 307668 164336
rect 274140 164296 274146 164308
rect 307662 164296 307668 164308
rect 307720 164296 307726 164348
rect 258810 164228 258816 164280
rect 258868 164268 258874 164280
rect 307294 164268 307300 164280
rect 258868 164240 307300 164268
rect 258868 164228 258874 164240
rect 307294 164228 307300 164240
rect 307352 164228 307358 164280
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 50338 164200 50344 164212
rect 3292 164172 50344 164200
rect 3292 164160 3298 164172
rect 50338 164160 50344 164172
rect 50396 164160 50402 164212
rect 166350 164160 166356 164212
rect 166408 164200 166414 164212
rect 214006 164200 214012 164212
rect 166408 164172 214012 164200
rect 166408 164160 166414 164172
rect 214006 164160 214012 164172
rect 214064 164160 214070 164212
rect 252462 164160 252468 164212
rect 252520 164200 252526 164212
rect 267734 164200 267740 164212
rect 252520 164172 267740 164200
rect 252520 164160 252526 164172
rect 267734 164160 267740 164172
rect 267792 164160 267798 164212
rect 324406 164160 324412 164212
rect 324464 164200 324470 164212
rect 345290 164200 345296 164212
rect 324464 164172 345296 164200
rect 324464 164160 324470 164172
rect 345290 164160 345296 164172
rect 345348 164160 345354 164212
rect 170674 164092 170680 164144
rect 170732 164132 170738 164144
rect 213914 164132 213920 164144
rect 170732 164104 213920 164132
rect 170732 164092 170738 164104
rect 213914 164092 213920 164104
rect 213972 164092 213978 164144
rect 251450 164092 251456 164144
rect 251508 164132 251514 164144
rect 253934 164132 253940 164144
rect 251508 164104 253940 164132
rect 251508 164092 251514 164104
rect 253934 164092 253940 164104
rect 253992 164092 253998 164144
rect 324314 164092 324320 164144
rect 324372 164132 324378 164144
rect 334066 164132 334072 164144
rect 324372 164104 334072 164132
rect 324372 164092 324378 164104
rect 334066 164092 334072 164104
rect 334124 164092 334130 164144
rect 297450 163004 297456 163056
rect 297508 163044 297514 163056
rect 307570 163044 307576 163056
rect 297508 163016 307576 163044
rect 297508 163004 297514 163016
rect 307570 163004 307576 163016
rect 307628 163004 307634 163056
rect 269758 162936 269764 162988
rect 269816 162976 269822 162988
rect 307478 162976 307484 162988
rect 269816 162948 307484 162976
rect 269816 162936 269822 162948
rect 307478 162936 307484 162948
rect 307536 162936 307542 162988
rect 261478 162868 261484 162920
rect 261536 162908 261542 162920
rect 307662 162908 307668 162920
rect 261536 162880 307668 162908
rect 261536 162868 261542 162880
rect 307662 162868 307668 162880
rect 307720 162868 307726 162920
rect 170398 162800 170404 162852
rect 170456 162840 170462 162852
rect 213914 162840 213920 162852
rect 170456 162812 213920 162840
rect 170456 162800 170462 162812
rect 213914 162800 213920 162812
rect 213972 162800 213978 162852
rect 252370 162800 252376 162852
rect 252428 162840 252434 162852
rect 266354 162840 266360 162852
rect 252428 162812 266360 162840
rect 252428 162800 252434 162812
rect 266354 162800 266360 162812
rect 266412 162800 266418 162852
rect 324314 162800 324320 162852
rect 324372 162840 324378 162852
rect 331490 162840 331496 162852
rect 324372 162812 331496 162840
rect 324372 162800 324378 162812
rect 331490 162800 331496 162812
rect 331548 162800 331554 162852
rect 252278 162732 252284 162784
rect 252336 162772 252342 162784
rect 263686 162772 263692 162784
rect 252336 162744 263692 162772
rect 252336 162732 252342 162744
rect 263686 162732 263692 162744
rect 263744 162732 263750 162784
rect 252462 162664 252468 162716
rect 252520 162704 252526 162716
rect 262398 162704 262404 162716
rect 252520 162676 262404 162704
rect 252520 162664 252526 162676
rect 262398 162664 262404 162676
rect 262456 162664 262462 162716
rect 324314 161848 324320 161900
rect 324372 161888 324378 161900
rect 327258 161888 327264 161900
rect 324372 161860 327264 161888
rect 324372 161848 324378 161860
rect 327258 161848 327264 161860
rect 327316 161848 327322 161900
rect 289354 161576 289360 161628
rect 289412 161616 289418 161628
rect 307570 161616 307576 161628
rect 289412 161588 307576 161616
rect 289412 161576 289418 161588
rect 307570 161576 307576 161588
rect 307628 161576 307634 161628
rect 286318 161508 286324 161560
rect 286376 161548 286382 161560
rect 307662 161548 307668 161560
rect 286376 161520 307668 161548
rect 286376 161508 286382 161520
rect 307662 161508 307668 161520
rect 307720 161508 307726 161560
rect 253198 161440 253204 161492
rect 253256 161480 253262 161492
rect 307478 161480 307484 161492
rect 253256 161452 307484 161480
rect 253256 161440 253262 161452
rect 307478 161440 307484 161452
rect 307536 161440 307542 161492
rect 171778 161372 171784 161424
rect 171836 161412 171842 161424
rect 214006 161412 214012 161424
rect 171836 161384 214012 161412
rect 171836 161372 171842 161384
rect 214006 161372 214012 161384
rect 214064 161372 214070 161424
rect 324314 161372 324320 161424
rect 324372 161412 324378 161424
rect 345106 161412 345112 161424
rect 324372 161384 345112 161412
rect 324372 161372 324378 161384
rect 345106 161372 345112 161384
rect 345164 161372 345170 161424
rect 195330 161304 195336 161356
rect 195388 161344 195394 161356
rect 213914 161344 213920 161356
rect 195388 161316 213920 161344
rect 195388 161304 195394 161316
rect 213914 161304 213920 161316
rect 213972 161304 213978 161356
rect 324406 161304 324412 161356
rect 324464 161344 324470 161356
rect 338390 161344 338396 161356
rect 324464 161316 338396 161344
rect 324464 161304 324470 161316
rect 338390 161304 338396 161316
rect 338448 161304 338454 161356
rect 252462 160760 252468 160812
rect 252520 160800 252526 160812
rect 259730 160800 259736 160812
rect 252520 160772 259736 160800
rect 252520 160760 252526 160772
rect 259730 160760 259736 160772
rect 259788 160760 259794 160812
rect 267274 160692 267280 160744
rect 267332 160732 267338 160744
rect 307294 160732 307300 160744
rect 267332 160704 307300 160732
rect 267332 160692 267338 160704
rect 307294 160692 307300 160704
rect 307352 160692 307358 160744
rect 304534 160148 304540 160200
rect 304592 160188 304598 160200
rect 307662 160188 307668 160200
rect 304592 160160 307668 160188
rect 304592 160148 304598 160160
rect 307662 160148 307668 160160
rect 307720 160148 307726 160200
rect 260098 160080 260104 160132
rect 260156 160120 260162 160132
rect 307570 160120 307576 160132
rect 260156 160092 307576 160120
rect 260156 160080 260162 160092
rect 307570 160080 307576 160092
rect 307628 160080 307634 160132
rect 173158 160012 173164 160064
rect 173216 160052 173222 160064
rect 213914 160052 213920 160064
rect 173216 160024 213920 160052
rect 173216 160012 173222 160024
rect 213914 160012 213920 160024
rect 213972 160012 213978 160064
rect 252462 160012 252468 160064
rect 252520 160052 252526 160064
rect 267826 160052 267832 160064
rect 252520 160024 267832 160052
rect 252520 160012 252526 160024
rect 267826 160012 267832 160024
rect 267884 160012 267890 160064
rect 324314 160012 324320 160064
rect 324372 160052 324378 160064
rect 345198 160052 345204 160064
rect 324372 160024 345204 160052
rect 324372 160012 324378 160024
rect 345198 160012 345204 160024
rect 345256 160012 345262 160064
rect 252002 159944 252008 159996
rect 252060 159984 252066 159996
rect 255314 159984 255320 159996
rect 252060 159956 255320 159984
rect 252060 159944 252066 159956
rect 255314 159944 255320 159956
rect 255372 159944 255378 159996
rect 298738 158856 298744 158908
rect 298796 158896 298802 158908
rect 306558 158896 306564 158908
rect 298796 158868 306564 158896
rect 298796 158856 298802 158868
rect 306558 158856 306564 158868
rect 306616 158856 306622 158908
rect 262950 158788 262956 158840
rect 263008 158828 263014 158840
rect 307294 158828 307300 158840
rect 263008 158800 307300 158828
rect 263008 158788 263014 158800
rect 307294 158788 307300 158800
rect 307352 158788 307358 158840
rect 258718 158720 258724 158772
rect 258776 158760 258782 158772
rect 307662 158760 307668 158772
rect 258776 158732 307668 158760
rect 258776 158720 258782 158732
rect 307662 158720 307668 158732
rect 307720 158720 307726 158772
rect 167638 158652 167644 158704
rect 167696 158692 167702 158704
rect 213914 158692 213920 158704
rect 167696 158664 213920 158692
rect 167696 158652 167702 158664
rect 213914 158652 213920 158664
rect 213972 158652 213978 158704
rect 324406 158652 324412 158704
rect 324464 158692 324470 158704
rect 341150 158692 341156 158704
rect 324464 158664 341156 158692
rect 324464 158652 324470 158664
rect 341150 158652 341156 158664
rect 341208 158652 341214 158704
rect 186958 158584 186964 158636
rect 187016 158624 187022 158636
rect 214006 158624 214012 158636
rect 187016 158596 214012 158624
rect 187016 158584 187022 158596
rect 214006 158584 214012 158596
rect 214064 158584 214070 158636
rect 324314 158584 324320 158636
rect 324372 158624 324378 158636
rect 336918 158624 336924 158636
rect 324372 158596 336924 158624
rect 324372 158584 324378 158596
rect 336918 158584 336924 158596
rect 336976 158584 336982 158636
rect 256142 157564 256148 157616
rect 256200 157604 256206 157616
rect 306926 157604 306932 157616
rect 256200 157576 306932 157604
rect 256200 157564 256206 157576
rect 306926 157564 306932 157576
rect 306984 157564 306990 157616
rect 295978 157496 295984 157548
rect 296036 157536 296042 157548
rect 307662 157536 307668 157548
rect 296036 157508 307668 157536
rect 296036 157496 296042 157508
rect 307662 157496 307668 157508
rect 307720 157496 307726 157548
rect 267090 157428 267096 157480
rect 267148 157468 267154 157480
rect 307570 157468 307576 157480
rect 267148 157440 307576 157468
rect 267148 157428 267154 157440
rect 307570 157428 307576 157440
rect 307628 157428 307634 157480
rect 169018 157292 169024 157344
rect 169076 157332 169082 157344
rect 214006 157332 214012 157344
rect 169076 157304 214012 157332
rect 169076 157292 169082 157304
rect 214006 157292 214012 157304
rect 214064 157292 214070 157344
rect 252462 157292 252468 157344
rect 252520 157332 252526 157344
rect 281534 157332 281540 157344
rect 252520 157304 281540 157332
rect 252520 157292 252526 157304
rect 281534 157292 281540 157304
rect 281592 157292 281598 157344
rect 324314 157292 324320 157344
rect 324372 157332 324378 157344
rect 328638 157332 328644 157344
rect 324372 157304 328644 157332
rect 324372 157292 324378 157304
rect 328638 157292 328644 157304
rect 328696 157292 328702 157344
rect 209038 157224 209044 157276
rect 209096 157264 209102 157276
rect 213914 157264 213920 157276
rect 209096 157236 213920 157264
rect 209096 157224 209102 157236
rect 213914 157224 213920 157236
rect 213972 157224 213978 157276
rect 252370 157224 252376 157276
rect 252428 157264 252434 157276
rect 270678 157264 270684 157276
rect 252428 157236 270684 157264
rect 252428 157224 252434 157236
rect 270678 157224 270684 157236
rect 270736 157224 270742 157276
rect 252462 157156 252468 157208
rect 252520 157196 252526 157208
rect 263778 157196 263784 157208
rect 252520 157168 263784 157196
rect 252520 157156 252526 157168
rect 263778 157156 263784 157168
rect 263836 157156 263842 157208
rect 296162 156068 296168 156120
rect 296220 156108 296226 156120
rect 307662 156108 307668 156120
rect 296220 156080 307668 156108
rect 296220 156068 296226 156080
rect 307662 156068 307668 156080
rect 307720 156068 307726 156120
rect 262858 156000 262864 156052
rect 262916 156040 262922 156052
rect 307478 156040 307484 156052
rect 262916 156012 307484 156040
rect 262916 156000 262922 156012
rect 307478 156000 307484 156012
rect 307536 156000 307542 156052
rect 260190 155932 260196 155984
rect 260248 155972 260254 155984
rect 307570 155972 307576 155984
rect 260248 155944 307576 155972
rect 260248 155932 260254 155944
rect 307570 155932 307576 155944
rect 307628 155932 307634 155984
rect 169202 155864 169208 155916
rect 169260 155904 169266 155916
rect 213914 155904 213920 155916
rect 169260 155876 213920 155904
rect 169260 155864 169266 155876
rect 213914 155864 213920 155876
rect 213972 155864 213978 155916
rect 252370 155864 252376 155916
rect 252428 155904 252434 155916
rect 265066 155904 265072 155916
rect 252428 155876 265072 155904
rect 252428 155864 252434 155876
rect 265066 155864 265072 155876
rect 265124 155864 265130 155916
rect 324406 155864 324412 155916
rect 324464 155904 324470 155916
rect 347958 155904 347964 155916
rect 324464 155876 347964 155904
rect 324464 155864 324470 155876
rect 347958 155864 347964 155876
rect 348016 155864 348022 155916
rect 252462 155796 252468 155848
rect 252520 155836 252526 155848
rect 261110 155836 261116 155848
rect 252520 155808 261116 155836
rect 252520 155796 252526 155808
rect 261110 155796 261116 155808
rect 261168 155796 261174 155848
rect 324314 155796 324320 155848
rect 324372 155836 324378 155848
rect 346486 155836 346492 155848
rect 324372 155808 346492 155836
rect 324372 155796 324378 155808
rect 346486 155796 346492 155808
rect 346544 155796 346550 155848
rect 251450 155728 251456 155780
rect 251508 155768 251514 155780
rect 254118 155768 254124 155780
rect 251508 155740 254124 155768
rect 251508 155728 251514 155740
rect 254118 155728 254124 155740
rect 254176 155728 254182 155780
rect 300210 154708 300216 154760
rect 300268 154748 300274 154760
rect 307662 154748 307668 154760
rect 300268 154720 307668 154748
rect 300268 154708 300274 154720
rect 307662 154708 307668 154720
rect 307720 154708 307726 154760
rect 285030 154640 285036 154692
rect 285088 154680 285094 154692
rect 306558 154680 306564 154692
rect 285088 154652 306564 154680
rect 285088 154640 285094 154652
rect 306558 154640 306564 154652
rect 306616 154640 306622 154692
rect 264514 154572 264520 154624
rect 264572 154612 264578 154624
rect 307294 154612 307300 154624
rect 264572 154584 307300 154612
rect 264572 154572 264578 154584
rect 307294 154572 307300 154584
rect 307352 154572 307358 154624
rect 252370 154504 252376 154556
rect 252428 154544 252434 154556
rect 271966 154544 271972 154556
rect 252428 154516 271972 154544
rect 252428 154504 252434 154516
rect 271966 154504 271972 154516
rect 272024 154504 272030 154556
rect 324314 154504 324320 154556
rect 324372 154544 324378 154556
rect 347866 154544 347872 154556
rect 324372 154516 347872 154544
rect 324372 154504 324378 154516
rect 347866 154504 347872 154516
rect 347924 154504 347930 154556
rect 252462 154436 252468 154488
rect 252520 154476 252526 154488
rect 267918 154476 267924 154488
rect 252520 154448 267924 154476
rect 252520 154436 252526 154448
rect 267918 154436 267924 154448
rect 267976 154436 267982 154488
rect 252278 154368 252284 154420
rect 252336 154408 252342 154420
rect 255498 154408 255504 154420
rect 252336 154380 255504 154408
rect 252336 154368 252342 154380
rect 255498 154368 255504 154380
rect 255556 154368 255562 154420
rect 324314 153756 324320 153808
rect 324372 153796 324378 153808
rect 327350 153796 327356 153808
rect 324372 153768 327356 153796
rect 324372 153756 324378 153768
rect 327350 153756 327356 153768
rect 327408 153756 327414 153808
rect 197998 153280 198004 153332
rect 198056 153320 198062 153332
rect 214006 153320 214012 153332
rect 198056 153292 214012 153320
rect 198056 153280 198062 153292
rect 214006 153280 214012 153292
rect 214064 153280 214070 153332
rect 303522 153280 303528 153332
rect 303580 153320 303586 153332
rect 307662 153320 307668 153332
rect 303580 153292 307668 153320
rect 303580 153280 303586 153292
rect 307662 153280 307668 153292
rect 307720 153280 307726 153332
rect 178678 153212 178684 153264
rect 178736 153252 178742 153264
rect 213914 153252 213920 153264
rect 178736 153224 213920 153252
rect 178736 153212 178742 153224
rect 213914 153212 213920 153224
rect 213972 153212 213978 153264
rect 282454 153212 282460 153264
rect 282512 153252 282518 153264
rect 306558 153252 306564 153264
rect 282512 153224 306564 153252
rect 282512 153212 282518 153224
rect 306558 153212 306564 153224
rect 306616 153212 306622 153264
rect 324406 153144 324412 153196
rect 324464 153184 324470 153196
rect 342530 153184 342536 153196
rect 324464 153156 342536 153184
rect 324464 153144 324470 153156
rect 342530 153144 342536 153156
rect 342588 153144 342594 153196
rect 393958 153144 393964 153196
rect 394016 153184 394022 153196
rect 579798 153184 579804 153196
rect 394016 153156 579804 153184
rect 394016 153144 394022 153156
rect 579798 153144 579804 153156
rect 579856 153144 579862 153196
rect 252462 153076 252468 153128
rect 252520 153116 252526 153128
rect 269206 153116 269212 153128
rect 252520 153088 269212 153116
rect 252520 153076 252526 153088
rect 269206 153076 269212 153088
rect 269264 153076 269270 153128
rect 304258 151920 304264 151972
rect 304316 151960 304322 151972
rect 307570 151960 307576 151972
rect 304316 151932 307576 151960
rect 304316 151920 304322 151932
rect 307570 151920 307576 151932
rect 307628 151920 307634 151972
rect 268470 151852 268476 151904
rect 268528 151892 268534 151904
rect 307662 151892 307668 151904
rect 268528 151864 307668 151892
rect 268528 151852 268534 151864
rect 307662 151852 307668 151864
rect 307720 151852 307726 151904
rect 177574 151784 177580 151836
rect 177632 151824 177638 151836
rect 213914 151824 213920 151836
rect 177632 151796 213920 151824
rect 177632 151784 177638 151796
rect 213914 151784 213920 151796
rect 213972 151784 213978 151836
rect 256050 151784 256056 151836
rect 256108 151824 256114 151836
rect 307478 151824 307484 151836
rect 256108 151796 307484 151824
rect 256108 151784 256114 151796
rect 307478 151784 307484 151796
rect 307536 151784 307542 151836
rect 252462 151716 252468 151768
rect 252520 151756 252526 151768
rect 276014 151756 276020 151768
rect 252520 151728 276020 151756
rect 252520 151716 252526 151728
rect 276014 151716 276020 151728
rect 276072 151716 276078 151768
rect 324314 151648 324320 151700
rect 324372 151688 324378 151700
rect 347774 151688 347780 151700
rect 324372 151660 347780 151688
rect 324372 151648 324378 151660
rect 347774 151648 347780 151660
rect 347832 151648 347838 151700
rect 252002 151444 252008 151496
rect 252060 151484 252066 151496
rect 254210 151484 254216 151496
rect 252060 151456 254216 151484
rect 252060 151444 252066 151456
rect 254210 151444 254216 151456
rect 254268 151444 254274 151496
rect 173250 151036 173256 151088
rect 173308 151076 173314 151088
rect 214374 151076 214380 151088
rect 173308 151048 214380 151076
rect 173308 151036 173314 151048
rect 214374 151036 214380 151048
rect 214432 151036 214438 151088
rect 287974 150560 287980 150612
rect 288032 150600 288038 150612
rect 307662 150600 307668 150612
rect 288032 150572 307668 150600
rect 288032 150560 288038 150572
rect 307662 150560 307668 150572
rect 307720 150560 307726 150612
rect 264330 150492 264336 150544
rect 264388 150532 264394 150544
rect 307294 150532 307300 150544
rect 264388 150504 307300 150532
rect 264388 150492 264394 150504
rect 307294 150492 307300 150504
rect 307352 150492 307358 150544
rect 175918 150424 175924 150476
rect 175976 150464 175982 150476
rect 214006 150464 214012 150476
rect 175976 150436 214012 150464
rect 175976 150424 175982 150436
rect 214006 150424 214012 150436
rect 214064 150424 214070 150476
rect 254578 150424 254584 150476
rect 254636 150464 254642 150476
rect 306926 150464 306932 150476
rect 254636 150436 306932 150464
rect 254636 150424 254642 150436
rect 306926 150424 306932 150436
rect 306984 150424 306990 150476
rect 3510 150356 3516 150408
rect 3568 150396 3574 150408
rect 25498 150396 25504 150408
rect 3568 150368 25504 150396
rect 3568 150356 3574 150368
rect 25498 150356 25504 150368
rect 25556 150356 25562 150408
rect 169110 150356 169116 150408
rect 169168 150396 169174 150408
rect 213914 150396 213920 150408
rect 169168 150368 213920 150396
rect 169168 150356 169174 150368
rect 213914 150356 213920 150368
rect 213972 150356 213978 150408
rect 252462 150356 252468 150408
rect 252520 150396 252526 150408
rect 278774 150396 278780 150408
rect 252520 150368 278780 150396
rect 252520 150356 252526 150368
rect 278774 150356 278780 150368
rect 278832 150356 278838 150408
rect 324314 150356 324320 150408
rect 324372 150396 324378 150408
rect 334250 150396 334256 150408
rect 324372 150368 334256 150396
rect 324372 150356 324378 150368
rect 334250 150356 334256 150368
rect 334308 150356 334314 150408
rect 252370 150288 252376 150340
rect 252428 150328 252434 150340
rect 273254 150328 273260 150340
rect 252428 150300 273260 150328
rect 252428 150288 252434 150300
rect 273254 150288 273260 150300
rect 273312 150288 273318 150340
rect 252278 150220 252284 150272
rect 252336 150260 252342 150272
rect 256786 150260 256792 150272
rect 252336 150232 256792 150260
rect 252336 150220 252342 150232
rect 256786 150220 256792 150232
rect 256844 150220 256850 150272
rect 324406 150220 324412 150272
rect 324464 150260 324470 150272
rect 327166 150260 327172 150272
rect 324464 150232 327172 150260
rect 324464 150220 324470 150232
rect 327166 150220 327172 150232
rect 327224 150220 327230 150272
rect 299106 149744 299112 149796
rect 299164 149784 299170 149796
rect 306650 149784 306656 149796
rect 299164 149756 306656 149784
rect 299164 149744 299170 149756
rect 306650 149744 306656 149756
rect 306708 149744 306714 149796
rect 257338 149676 257344 149728
rect 257396 149716 257402 149728
rect 307110 149716 307116 149728
rect 257396 149688 307116 149716
rect 257396 149676 257402 149688
rect 307110 149676 307116 149688
rect 307168 149676 307174 149728
rect 281074 149064 281080 149116
rect 281132 149104 281138 149116
rect 307662 149104 307668 149116
rect 281132 149076 307668 149104
rect 281132 149064 281138 149076
rect 307662 149064 307668 149076
rect 307720 149064 307726 149116
rect 166258 148996 166264 149048
rect 166316 149036 166322 149048
rect 213914 149036 213920 149048
rect 166316 149008 213920 149036
rect 166316 148996 166322 149008
rect 213914 148996 213920 149008
rect 213972 148996 213978 149048
rect 252462 148996 252468 149048
rect 252520 149036 252526 149048
rect 280154 149036 280160 149048
rect 252520 149008 280160 149036
rect 252520 148996 252526 149008
rect 280154 148996 280160 149008
rect 280212 148996 280218 149048
rect 324314 148996 324320 149048
rect 324372 149036 324378 149048
rect 343726 149036 343732 149048
rect 324372 149008 343732 149036
rect 324372 148996 324378 149008
rect 343726 148996 343732 149008
rect 343784 148996 343790 149048
rect 252370 148928 252376 148980
rect 252428 148968 252434 148980
rect 276106 148968 276112 148980
rect 252428 148940 276112 148968
rect 252428 148928 252434 148940
rect 276106 148928 276112 148940
rect 276164 148928 276170 148980
rect 264422 147772 264428 147824
rect 264480 147812 264486 147824
rect 306558 147812 306564 147824
rect 264480 147784 306564 147812
rect 264480 147772 264486 147784
rect 306558 147772 306564 147784
rect 306616 147772 306622 147824
rect 167730 147636 167736 147688
rect 167788 147676 167794 147688
rect 213914 147676 213920 147688
rect 167788 147648 213920 147676
rect 167788 147636 167794 147648
rect 213914 147636 213920 147648
rect 213972 147636 213978 147688
rect 301774 147636 301780 147688
rect 301832 147676 301838 147688
rect 307662 147676 307668 147688
rect 301832 147648 307668 147676
rect 301832 147636 301838 147648
rect 307662 147636 307668 147648
rect 307720 147636 307726 147688
rect 252462 147568 252468 147620
rect 252520 147608 252526 147620
rect 274726 147608 274732 147620
rect 252520 147580 274732 147608
rect 252520 147568 252526 147580
rect 274726 147568 274732 147580
rect 274784 147568 274790 147620
rect 324314 147568 324320 147620
rect 324372 147608 324378 147620
rect 335354 147608 335360 147620
rect 324372 147580 335360 147608
rect 324372 147568 324378 147580
rect 335354 147568 335360 147580
rect 335412 147568 335418 147620
rect 251266 147500 251272 147552
rect 251324 147540 251330 147552
rect 254026 147540 254032 147552
rect 251324 147512 254032 147540
rect 251324 147500 251330 147512
rect 254026 147500 254032 147512
rect 254084 147500 254090 147552
rect 290642 146888 290648 146940
rect 290700 146928 290706 146940
rect 307202 146928 307208 146940
rect 290700 146900 307208 146928
rect 290700 146888 290706 146900
rect 307202 146888 307208 146900
rect 307260 146888 307266 146940
rect 210418 146344 210424 146396
rect 210476 146384 210482 146396
rect 214006 146384 214012 146396
rect 210476 146356 214012 146384
rect 210476 146344 210482 146356
rect 214006 146344 214012 146356
rect 214064 146344 214070 146396
rect 255958 146344 255964 146396
rect 256016 146384 256022 146396
rect 307294 146384 307300 146396
rect 256016 146356 307300 146384
rect 256016 146344 256022 146356
rect 307294 146344 307300 146356
rect 307352 146344 307358 146396
rect 174538 146276 174544 146328
rect 174596 146316 174602 146328
rect 213914 146316 213920 146328
rect 174596 146288 213920 146316
rect 174596 146276 174602 146288
rect 213914 146276 213920 146288
rect 213972 146276 213978 146328
rect 254670 146276 254676 146328
rect 254728 146316 254734 146328
rect 306926 146316 306932 146328
rect 254728 146288 306932 146316
rect 254728 146276 254734 146288
rect 306926 146276 306932 146288
rect 306984 146276 306990 146328
rect 252278 146208 252284 146260
rect 252336 146248 252342 146260
rect 273346 146248 273352 146260
rect 252336 146220 273352 146248
rect 252336 146208 252342 146220
rect 273346 146208 273352 146220
rect 273404 146208 273410 146260
rect 324314 146208 324320 146260
rect 324372 146248 324378 146260
rect 339770 146248 339776 146260
rect 324372 146220 339776 146248
rect 324372 146208 324378 146220
rect 339770 146208 339776 146220
rect 339828 146208 339834 146260
rect 252462 146140 252468 146192
rect 252520 146180 252526 146192
rect 273438 146180 273444 146192
rect 252520 146152 273444 146180
rect 252520 146140 252526 146152
rect 273438 146140 273444 146152
rect 273496 146140 273502 146192
rect 324406 146140 324412 146192
rect 324464 146180 324470 146192
rect 328730 146180 328736 146192
rect 324464 146152 328736 146180
rect 324464 146140 324470 146152
rect 328730 146140 328736 146152
rect 328788 146140 328794 146192
rect 252370 146072 252376 146124
rect 252428 146112 252434 146124
rect 262306 146112 262312 146124
rect 252428 146084 262312 146112
rect 252428 146072 252434 146084
rect 262306 146072 262312 146084
rect 262364 146072 262370 146124
rect 292114 145596 292120 145648
rect 292172 145636 292178 145648
rect 307570 145636 307576 145648
rect 292172 145608 307576 145636
rect 292172 145596 292178 145608
rect 307570 145596 307576 145608
rect 307628 145596 307634 145648
rect 252002 145528 252008 145580
rect 252060 145568 252066 145580
rect 264238 145568 264244 145580
rect 252060 145540 264244 145568
rect 252060 145528 252066 145540
rect 264238 145528 264244 145540
rect 264296 145528 264302 145580
rect 285214 145528 285220 145580
rect 285272 145568 285278 145580
rect 307478 145568 307484 145580
rect 285272 145540 307484 145568
rect 285272 145528 285278 145540
rect 307478 145528 307484 145540
rect 307536 145528 307542 145580
rect 173158 144984 173164 145036
rect 173216 145024 173222 145036
rect 214006 145024 214012 145036
rect 173216 144996 214012 145024
rect 173216 144984 173222 144996
rect 214006 144984 214012 144996
rect 214064 144984 214070 145036
rect 169018 144916 169024 144968
rect 169076 144956 169082 144968
rect 213914 144956 213920 144968
rect 169076 144928 213920 144956
rect 169076 144916 169082 144928
rect 213914 144916 213920 144928
rect 213972 144916 213978 144968
rect 252462 144848 252468 144900
rect 252520 144888 252526 144900
rect 266446 144888 266452 144900
rect 252520 144860 266452 144888
rect 252520 144848 252526 144860
rect 266446 144848 266452 144860
rect 266504 144848 266510 144900
rect 324314 144848 324320 144900
rect 324372 144888 324378 144900
rect 331398 144888 331404 144900
rect 324372 144860 331404 144888
rect 324372 144848 324378 144860
rect 331398 144848 331404 144860
rect 331456 144848 331462 144900
rect 324406 144780 324412 144832
rect 324464 144820 324470 144832
rect 329926 144820 329932 144832
rect 324464 144792 329932 144820
rect 324464 144780 324470 144792
rect 329926 144780 329932 144792
rect 329984 144780 329990 144832
rect 299014 143692 299020 143744
rect 299072 143732 299078 143744
rect 307478 143732 307484 143744
rect 299072 143704 307484 143732
rect 299072 143692 299078 143704
rect 307478 143692 307484 143704
rect 307536 143692 307542 143744
rect 202138 143624 202144 143676
rect 202196 143664 202202 143676
rect 213914 143664 213920 143676
rect 202196 143636 213920 143664
rect 202196 143624 202202 143636
rect 213914 143624 213920 143636
rect 213972 143624 213978 143676
rect 268562 143624 268568 143676
rect 268620 143664 268626 143676
rect 307570 143664 307576 143676
rect 268620 143636 307576 143664
rect 268620 143624 268626 143636
rect 307570 143624 307576 143636
rect 307628 143624 307634 143676
rect 166258 143556 166264 143608
rect 166316 143596 166322 143608
rect 214006 143596 214012 143608
rect 166316 143568 214012 143596
rect 166316 143556 166322 143568
rect 214006 143556 214012 143568
rect 214064 143556 214070 143608
rect 253290 143556 253296 143608
rect 253348 143596 253354 143608
rect 307662 143596 307668 143608
rect 253348 143568 307668 143596
rect 253348 143556 253354 143568
rect 307662 143556 307668 143568
rect 307720 143556 307726 143608
rect 252370 143488 252376 143540
rect 252428 143528 252434 143540
rect 270494 143528 270500 143540
rect 252428 143500 270500 143528
rect 252428 143488 252434 143500
rect 270494 143488 270500 143500
rect 270552 143488 270558 143540
rect 324406 143488 324412 143540
rect 324464 143528 324470 143540
rect 351914 143528 351920 143540
rect 324464 143500 351920 143528
rect 324464 143488 324470 143500
rect 351914 143488 351920 143500
rect 351972 143488 351978 143540
rect 252462 143420 252468 143472
rect 252520 143460 252526 143472
rect 269114 143460 269120 143472
rect 252520 143432 269120 143460
rect 252520 143420 252526 143432
rect 269114 143420 269120 143432
rect 269172 143420 269178 143472
rect 324314 143420 324320 143472
rect 324372 143460 324378 143472
rect 334158 143460 334164 143472
rect 324372 143432 334164 143460
rect 324372 143420 324378 143432
rect 334158 143420 334164 143432
rect 334216 143420 334222 143472
rect 251910 142808 251916 142860
rect 251968 142848 251974 142860
rect 280798 142848 280804 142860
rect 251968 142820 280804 142848
rect 251968 142808 251974 142820
rect 280798 142808 280804 142820
rect 280856 142808 280862 142860
rect 300302 142264 300308 142316
rect 300360 142304 300366 142316
rect 307662 142304 307668 142316
rect 300360 142276 307668 142304
rect 300360 142264 300366 142276
rect 307662 142264 307668 142276
rect 307720 142264 307726 142316
rect 280982 142196 280988 142248
rect 281040 142236 281046 142248
rect 306558 142236 306564 142248
rect 281040 142208 306564 142236
rect 281040 142196 281046 142208
rect 306558 142196 306564 142208
rect 306616 142196 306622 142248
rect 206370 142128 206376 142180
rect 206428 142168 206434 142180
rect 213914 142168 213920 142180
rect 206428 142140 213920 142168
rect 206428 142128 206434 142140
rect 213914 142128 213920 142140
rect 213972 142128 213978 142180
rect 269942 142128 269948 142180
rect 270000 142168 270006 142180
rect 307570 142168 307576 142180
rect 270000 142140 307576 142168
rect 270000 142128 270006 142140
rect 307570 142128 307576 142140
rect 307628 142128 307634 142180
rect 252462 142060 252468 142112
rect 252520 142100 252526 142112
rect 262214 142100 262220 142112
rect 252520 142072 262220 142100
rect 252520 142060 252526 142072
rect 262214 142060 262220 142072
rect 262272 142060 262278 142112
rect 324406 142060 324412 142112
rect 324464 142100 324470 142112
rect 342254 142100 342260 142112
rect 324464 142072 342260 142100
rect 324464 142060 324470 142072
rect 342254 142060 342260 142072
rect 342312 142060 342318 142112
rect 324314 141992 324320 142044
rect 324372 142032 324378 142044
rect 339586 142032 339592 142044
rect 324372 142004 339592 142032
rect 324372 141992 324378 142004
rect 339586 141992 339592 142004
rect 339644 141992 339650 142044
rect 253382 141380 253388 141432
rect 253440 141420 253446 141432
rect 307478 141420 307484 141432
rect 253440 141392 307484 141420
rect 253440 141380 253446 141392
rect 307478 141380 307484 141392
rect 307536 141380 307542 141432
rect 275278 140904 275284 140956
rect 275336 140944 275342 140956
rect 307662 140944 307668 140956
rect 275336 140916 307668 140944
rect 275336 140904 275342 140916
rect 307662 140904 307668 140916
rect 307720 140904 307726 140956
rect 177390 140836 177396 140888
rect 177448 140876 177454 140888
rect 213914 140876 213920 140888
rect 177448 140848 213920 140876
rect 177448 140836 177454 140848
rect 213914 140836 213920 140848
rect 213972 140836 213978 140888
rect 294874 140836 294880 140888
rect 294932 140876 294938 140888
rect 306558 140876 306564 140888
rect 294932 140848 306564 140876
rect 294932 140836 294938 140848
rect 306558 140836 306564 140848
rect 306616 140836 306622 140888
rect 167638 140768 167644 140820
rect 167696 140808 167702 140820
rect 214006 140808 214012 140820
rect 167696 140780 214012 140808
rect 167696 140768 167702 140780
rect 214006 140768 214012 140780
rect 214064 140768 214070 140820
rect 304442 140768 304448 140820
rect 304500 140808 304506 140820
rect 307570 140808 307576 140820
rect 304500 140780 307576 140808
rect 304500 140768 304506 140780
rect 307570 140768 307576 140780
rect 307628 140768 307634 140820
rect 252462 140700 252468 140752
rect 252520 140740 252526 140752
rect 274634 140740 274640 140752
rect 252520 140712 274640 140740
rect 252520 140700 252526 140712
rect 274634 140700 274640 140712
rect 274692 140700 274698 140752
rect 324314 140700 324320 140752
rect 324372 140740 324378 140752
rect 329834 140740 329840 140752
rect 324372 140712 329840 140740
rect 324372 140700 324378 140712
rect 329834 140700 329840 140712
rect 329892 140700 329898 140752
rect 252370 140632 252376 140684
rect 252428 140672 252434 140684
rect 256970 140672 256976 140684
rect 252428 140644 256976 140672
rect 252428 140632 252434 140644
rect 256970 140632 256976 140644
rect 257028 140632 257034 140684
rect 257430 140020 257436 140072
rect 257488 140060 257494 140072
rect 307110 140060 307116 140072
rect 257488 140032 307116 140060
rect 257488 140020 257494 140032
rect 307110 140020 307116 140032
rect 307168 140020 307174 140072
rect 209038 139476 209044 139528
rect 209096 139516 209102 139528
rect 213914 139516 213920 139528
rect 209096 139488 213920 139516
rect 209096 139476 209102 139488
rect 213914 139476 213920 139488
rect 213972 139476 213978 139528
rect 289078 139476 289084 139528
rect 289136 139516 289142 139528
rect 306926 139516 306932 139528
rect 289136 139488 306932 139516
rect 289136 139476 289142 139488
rect 306926 139476 306932 139488
rect 306984 139476 306990 139528
rect 171778 139408 171784 139460
rect 171836 139448 171842 139460
rect 214006 139448 214012 139460
rect 171836 139420 214012 139448
rect 171836 139408 171842 139420
rect 214006 139408 214012 139420
rect 214064 139408 214070 139460
rect 279510 139408 279516 139460
rect 279568 139448 279574 139460
rect 307294 139448 307300 139460
rect 279568 139420 307300 139448
rect 279568 139408 279574 139420
rect 307294 139408 307300 139420
rect 307352 139408 307358 139460
rect 252278 139340 252284 139392
rect 252336 139380 252342 139392
rect 255590 139380 255596 139392
rect 252336 139352 255596 139380
rect 252336 139340 252342 139352
rect 255590 139340 255596 139352
rect 255648 139340 255654 139392
rect 324406 139340 324412 139392
rect 324464 139380 324470 139392
rect 332870 139380 332876 139392
rect 324464 139352 332876 139380
rect 324464 139340 324470 139352
rect 332870 139340 332876 139352
rect 332928 139340 332934 139392
rect 324314 139272 324320 139324
rect 324372 139312 324378 139324
rect 331306 139312 331312 139324
rect 324372 139284 331312 139312
rect 324372 139272 324378 139284
rect 331306 139272 331312 139284
rect 331364 139272 331370 139324
rect 252186 138660 252192 138712
rect 252244 138700 252250 138712
rect 265802 138700 265808 138712
rect 252244 138672 265808 138700
rect 252244 138660 252250 138672
rect 265802 138660 265808 138672
rect 265860 138660 265866 138712
rect 280798 138116 280804 138168
rect 280856 138156 280862 138168
rect 307662 138156 307668 138168
rect 280856 138128 307668 138156
rect 280856 138116 280862 138128
rect 307662 138116 307668 138128
rect 307720 138116 307726 138168
rect 266998 138048 267004 138100
rect 267056 138088 267062 138100
rect 307570 138088 307576 138100
rect 267056 138060 307576 138088
rect 267056 138048 267062 138060
rect 307570 138048 307576 138060
rect 307628 138048 307634 138100
rect 170398 137980 170404 138032
rect 170456 138020 170462 138032
rect 213914 138020 213920 138032
rect 170456 137992 213920 138020
rect 170456 137980 170462 137992
rect 213914 137980 213920 137992
rect 213972 137980 213978 138032
rect 250438 137980 250444 138032
rect 250496 138020 250502 138032
rect 306558 138020 306564 138032
rect 250496 137992 306564 138020
rect 250496 137980 250502 137992
rect 306558 137980 306564 137992
rect 306616 137980 306622 138032
rect 3510 137912 3516 137964
rect 3568 137952 3574 137964
rect 14458 137952 14464 137964
rect 3568 137924 14464 137952
rect 3568 137912 3574 137924
rect 14458 137912 14464 137924
rect 14516 137912 14522 137964
rect 252278 137912 252284 137964
rect 252336 137952 252342 137964
rect 277486 137952 277492 137964
rect 252336 137924 277492 137952
rect 252336 137912 252342 137924
rect 277486 137912 277492 137924
rect 277544 137912 277550 137964
rect 324314 137912 324320 137964
rect 324372 137952 324378 137964
rect 343634 137952 343640 137964
rect 324372 137924 343640 137952
rect 324372 137912 324378 137924
rect 343634 137912 343640 137924
rect 343692 137912 343698 137964
rect 252370 137844 252376 137896
rect 252428 137884 252434 137896
rect 277394 137884 277400 137896
rect 252428 137856 277400 137884
rect 252428 137844 252434 137856
rect 277394 137844 277400 137856
rect 277452 137844 277458 137896
rect 324406 137844 324412 137896
rect 324464 137884 324470 137896
rect 335446 137884 335452 137896
rect 324464 137856 335452 137884
rect 324464 137844 324470 137856
rect 335446 137844 335452 137856
rect 335504 137844 335510 137896
rect 252462 137776 252468 137828
rect 252520 137816 252526 137828
rect 271874 137816 271880 137828
rect 252520 137788 271880 137816
rect 252520 137776 252526 137788
rect 271874 137776 271880 137788
rect 271932 137776 271938 137828
rect 251818 137300 251824 137352
rect 251876 137340 251882 137352
rect 295978 137340 295984 137352
rect 251876 137312 295984 137340
rect 251876 137300 251882 137312
rect 295978 137300 295984 137312
rect 296036 137300 296042 137352
rect 171962 137232 171968 137284
rect 172020 137272 172026 137284
rect 214558 137272 214564 137284
rect 172020 137244 214564 137272
rect 172020 137232 172026 137244
rect 214558 137232 214564 137244
rect 214616 137232 214622 137284
rect 253474 137232 253480 137284
rect 253532 137272 253538 137284
rect 307018 137272 307024 137284
rect 253532 137244 307024 137272
rect 253532 137232 253538 137244
rect 307018 137232 307024 137244
rect 307076 137232 307082 137284
rect 297358 136688 297364 136740
rect 297416 136728 297422 136740
rect 307662 136728 307668 136740
rect 297416 136700 307668 136728
rect 297416 136688 297422 136700
rect 307662 136688 307668 136700
rect 307720 136688 307726 136740
rect 204898 136620 204904 136672
rect 204956 136660 204962 136672
rect 213914 136660 213920 136672
rect 204956 136632 213920 136660
rect 204956 136620 204962 136632
rect 213914 136620 213920 136632
rect 213972 136620 213978 136672
rect 293218 136620 293224 136672
rect 293276 136660 293282 136672
rect 307570 136660 307576 136672
rect 293276 136632 307576 136660
rect 293276 136620 293282 136632
rect 307570 136620 307576 136632
rect 307628 136620 307634 136672
rect 252278 136552 252284 136604
rect 252336 136592 252342 136604
rect 287790 136592 287796 136604
rect 252336 136564 287796 136592
rect 252336 136552 252342 136564
rect 287790 136552 287796 136564
rect 287848 136552 287854 136604
rect 324314 136552 324320 136604
rect 324372 136592 324378 136604
rect 341058 136592 341064 136604
rect 324372 136564 341064 136592
rect 324372 136552 324378 136564
rect 341058 136552 341064 136564
rect 341116 136552 341122 136604
rect 252462 136484 252468 136536
rect 252520 136524 252526 136536
rect 270586 136524 270592 136536
rect 252520 136496 270592 136524
rect 252520 136484 252526 136496
rect 270586 136484 270592 136496
rect 270644 136484 270650 136536
rect 252370 136416 252376 136468
rect 252428 136456 252434 136468
rect 268378 136456 268384 136468
rect 252428 136428 268384 136456
rect 252428 136416 252434 136428
rect 268378 136416 268384 136428
rect 268436 136416 268442 136468
rect 324958 136212 324964 136264
rect 325016 136252 325022 136264
rect 327074 136252 327080 136264
rect 325016 136224 327080 136252
rect 325016 136212 325022 136224
rect 327074 136212 327080 136224
rect 327132 136212 327138 136264
rect 302878 135464 302884 135516
rect 302936 135504 302942 135516
rect 307294 135504 307300 135516
rect 302936 135476 307300 135504
rect 302936 135464 302942 135476
rect 307294 135464 307300 135476
rect 307352 135464 307358 135516
rect 287698 135396 287704 135448
rect 287756 135436 287762 135448
rect 306558 135436 306564 135448
rect 287756 135408 306564 135436
rect 287756 135396 287762 135408
rect 306558 135396 306564 135408
rect 306616 135396 306622 135448
rect 195238 135328 195244 135380
rect 195296 135368 195302 135380
rect 214006 135368 214012 135380
rect 195296 135340 214012 135368
rect 195296 135328 195302 135340
rect 214006 135328 214012 135340
rect 214064 135328 214070 135380
rect 283558 135328 283564 135380
rect 283616 135368 283622 135380
rect 307478 135368 307484 135380
rect 283616 135340 307484 135368
rect 283616 135328 283622 135340
rect 307478 135328 307484 135340
rect 307536 135328 307542 135380
rect 170490 135260 170496 135312
rect 170548 135300 170554 135312
rect 213914 135300 213920 135312
rect 170548 135272 213920 135300
rect 170548 135260 170554 135272
rect 213914 135260 213920 135272
rect 213972 135260 213978 135312
rect 278130 135260 278136 135312
rect 278188 135300 278194 135312
rect 307662 135300 307668 135312
rect 278188 135272 307668 135300
rect 278188 135260 278194 135272
rect 307662 135260 307668 135272
rect 307720 135260 307726 135312
rect 252462 135192 252468 135244
rect 252520 135232 252526 135244
rect 276658 135232 276664 135244
rect 252520 135204 276664 135232
rect 252520 135192 252526 135204
rect 276658 135192 276664 135204
rect 276716 135192 276722 135244
rect 307202 135192 307208 135244
rect 307260 135232 307266 135244
rect 307478 135232 307484 135244
rect 307260 135204 307484 135232
rect 307260 135192 307266 135204
rect 307478 135192 307484 135204
rect 307536 135192 307542 135244
rect 252370 135124 252376 135176
rect 252428 135164 252434 135176
rect 267182 135164 267188 135176
rect 252428 135136 267188 135164
rect 252428 135124 252434 135136
rect 267182 135124 267188 135136
rect 267240 135124 267246 135176
rect 324314 135124 324320 135176
rect 324372 135164 324378 135176
rect 339494 135164 339500 135176
rect 324372 135136 339500 135164
rect 324372 135124 324378 135136
rect 339494 135124 339500 135136
rect 339552 135124 339558 135176
rect 177482 133968 177488 134020
rect 177540 134008 177546 134020
rect 213914 134008 213920 134020
rect 177540 133980 213920 134008
rect 177540 133968 177546 133980
rect 213914 133968 213920 133980
rect 213972 133968 213978 134020
rect 291930 133968 291936 134020
rect 291988 134008 291994 134020
rect 307570 134008 307576 134020
rect 291988 133980 307576 134008
rect 291988 133968 291994 133980
rect 307570 133968 307576 133980
rect 307628 133968 307634 134020
rect 167822 133900 167828 133952
rect 167880 133940 167886 133952
rect 214006 133940 214012 133952
rect 167880 133912 214012 133940
rect 167880 133900 167886 133912
rect 214006 133900 214012 133912
rect 214064 133900 214070 133952
rect 276750 133900 276756 133952
rect 276808 133940 276814 133952
rect 307662 133940 307668 133952
rect 276808 133912 307668 133940
rect 276808 133900 276814 133912
rect 307662 133900 307668 133912
rect 307720 133900 307726 133952
rect 252370 133832 252376 133884
rect 252428 133872 252434 133884
rect 289170 133872 289176 133884
rect 252428 133844 289176 133872
rect 252428 133832 252434 133844
rect 289170 133832 289176 133844
rect 289228 133832 289234 133884
rect 324314 133832 324320 133884
rect 324372 133872 324378 133884
rect 330018 133872 330024 133884
rect 324372 133844 330024 133872
rect 324372 133832 324378 133844
rect 330018 133832 330024 133844
rect 330076 133832 330082 133884
rect 252462 133764 252468 133816
rect 252520 133804 252526 133816
rect 284938 133804 284944 133816
rect 252520 133776 284944 133804
rect 252520 133764 252526 133776
rect 284938 133764 284944 133776
rect 284996 133764 285002 133816
rect 286594 133152 286600 133204
rect 286652 133192 286658 133204
rect 306742 133192 306748 133204
rect 286652 133164 306748 133192
rect 286652 133152 286658 133164
rect 306742 133152 306748 133164
rect 306800 133152 306806 133204
rect 196710 132540 196716 132592
rect 196768 132580 196774 132592
rect 214006 132580 214012 132592
rect 196768 132552 214012 132580
rect 196768 132540 196774 132552
rect 214006 132540 214012 132552
rect 214064 132540 214070 132592
rect 290550 132540 290556 132592
rect 290608 132580 290614 132592
rect 307662 132580 307668 132592
rect 290608 132552 307668 132580
rect 290608 132540 290614 132552
rect 307662 132540 307668 132552
rect 307720 132540 307726 132592
rect 173342 132472 173348 132524
rect 173400 132512 173406 132524
rect 213914 132512 213920 132524
rect 173400 132484 213920 132512
rect 173400 132472 173406 132484
rect 213914 132472 213920 132484
rect 213972 132472 213978 132524
rect 282178 132472 282184 132524
rect 282236 132512 282242 132524
rect 307570 132512 307576 132524
rect 282236 132484 307576 132512
rect 282236 132472 282242 132484
rect 307570 132472 307576 132484
rect 307628 132472 307634 132524
rect 252278 132404 252284 132456
rect 252336 132444 252342 132456
rect 286410 132444 286416 132456
rect 252336 132416 286416 132444
rect 252336 132404 252342 132416
rect 286410 132404 286416 132416
rect 286468 132404 286474 132456
rect 324406 132404 324412 132456
rect 324464 132444 324470 132456
rect 346394 132444 346400 132456
rect 324464 132416 346400 132444
rect 324464 132404 324470 132416
rect 346394 132404 346400 132416
rect 346452 132404 346458 132456
rect 252462 132336 252468 132388
rect 252520 132376 252526 132388
rect 265710 132376 265716 132388
rect 252520 132348 265716 132376
rect 252520 132336 252526 132348
rect 265710 132336 265716 132348
rect 265768 132336 265774 132388
rect 324314 132336 324320 132388
rect 324372 132376 324378 132388
rect 345014 132376 345020 132388
rect 324372 132348 345020 132376
rect 324372 132336 324378 132348
rect 345014 132336 345020 132348
rect 345072 132336 345078 132388
rect 252370 131520 252376 131572
rect 252428 131560 252434 131572
rect 260282 131560 260288 131572
rect 252428 131532 260288 131560
rect 252428 131520 252434 131532
rect 260282 131520 260288 131532
rect 260340 131520 260346 131572
rect 294782 131248 294788 131300
rect 294840 131288 294846 131300
rect 307662 131288 307668 131300
rect 294840 131260 307668 131288
rect 294840 131248 294846 131260
rect 307662 131248 307668 131260
rect 307720 131248 307726 131300
rect 207658 131180 207664 131232
rect 207716 131220 207722 131232
rect 213914 131220 213920 131232
rect 207716 131192 213920 131220
rect 207716 131180 207722 131192
rect 213914 131180 213920 131192
rect 213972 131180 213978 131232
rect 278038 131180 278044 131232
rect 278096 131220 278102 131232
rect 307386 131220 307392 131232
rect 278096 131192 307392 131220
rect 278096 131180 278102 131192
rect 307386 131180 307392 131192
rect 307444 131180 307450 131232
rect 189718 131112 189724 131164
rect 189776 131152 189782 131164
rect 214006 131152 214012 131164
rect 189776 131124 214012 131152
rect 189776 131112 189782 131124
rect 214006 131112 214012 131124
rect 214064 131112 214070 131164
rect 271138 131112 271144 131164
rect 271196 131152 271202 131164
rect 307570 131152 307576 131164
rect 271196 131124 307576 131152
rect 271196 131112 271202 131124
rect 307570 131112 307576 131124
rect 307628 131112 307634 131164
rect 252278 131044 252284 131096
rect 252336 131084 252342 131096
rect 291838 131084 291844 131096
rect 252336 131056 291844 131084
rect 252336 131044 252342 131056
rect 291838 131044 291844 131056
rect 291896 131044 291902 131096
rect 324406 131044 324412 131096
rect 324464 131084 324470 131096
rect 342438 131084 342444 131096
rect 324464 131056 342444 131084
rect 324464 131044 324470 131056
rect 342438 131044 342444 131056
rect 342496 131044 342502 131096
rect 252462 130976 252468 131028
rect 252520 131016 252526 131028
rect 267274 131016 267280 131028
rect 252520 130988 267280 131016
rect 252520 130976 252526 130988
rect 267274 130976 267280 130988
rect 267332 130976 267338 131028
rect 324314 130976 324320 131028
rect 324372 131016 324378 131028
rect 331214 131016 331220 131028
rect 324372 130988 331220 131016
rect 324372 130976 324378 130988
rect 331214 130976 331220 130988
rect 331272 130976 331278 131028
rect 252370 130364 252376 130416
rect 252428 130404 252434 130416
rect 261570 130404 261576 130416
rect 252428 130376 261576 130404
rect 252428 130364 252434 130376
rect 261570 130364 261576 130376
rect 261628 130364 261634 130416
rect 296254 129888 296260 129940
rect 296312 129928 296318 129940
rect 307662 129928 307668 129940
rect 296312 129900 307668 129928
rect 296312 129888 296318 129900
rect 307662 129888 307668 129900
rect 307720 129888 307726 129940
rect 199378 129820 199384 129872
rect 199436 129860 199442 129872
rect 214006 129860 214012 129872
rect 199436 129832 214012 129860
rect 199436 129820 199442 129832
rect 214006 129820 214012 129832
rect 214064 129820 214070 129872
rect 285122 129820 285128 129872
rect 285180 129860 285186 129872
rect 307478 129860 307484 129872
rect 285180 129832 307484 129860
rect 285180 129820 285186 129832
rect 307478 129820 307484 129832
rect 307536 129820 307542 129872
rect 171870 129752 171876 129804
rect 171928 129792 171934 129804
rect 213914 129792 213920 129804
rect 171928 129764 213920 129792
rect 171928 129752 171934 129764
rect 213914 129752 213920 129764
rect 213972 129752 213978 129804
rect 273990 129752 273996 129804
rect 274048 129792 274054 129804
rect 307570 129792 307576 129804
rect 274048 129764 307576 129792
rect 274048 129752 274054 129764
rect 307570 129752 307576 129764
rect 307628 129752 307634 129804
rect 252462 129684 252468 129736
rect 252520 129724 252526 129736
rect 269850 129724 269856 129736
rect 252520 129696 269856 129724
rect 252520 129684 252526 129696
rect 269850 129684 269856 129696
rect 269908 129684 269914 129736
rect 324406 129684 324412 129736
rect 324464 129724 324470 129736
rect 346578 129724 346584 129736
rect 324464 129696 346584 129724
rect 324464 129684 324470 129696
rect 346578 129684 346584 129696
rect 346636 129684 346642 129736
rect 252278 129616 252284 129668
rect 252336 129656 252342 129668
rect 261662 129656 261668 129668
rect 252336 129628 261668 129656
rect 252336 129616 252342 129628
rect 261662 129616 261668 129628
rect 261720 129616 261726 129668
rect 324314 129616 324320 129668
rect 324372 129656 324378 129668
rect 330110 129656 330116 129668
rect 324372 129628 330116 129656
rect 324372 129616 324378 129628
rect 330110 129616 330116 129628
rect 330168 129616 330174 129668
rect 252002 129004 252008 129056
rect 252060 129044 252066 129056
rect 305730 129044 305736 129056
rect 252060 129016 305736 129044
rect 252060 129004 252066 129016
rect 305730 129004 305736 129016
rect 305788 129004 305794 129056
rect 301590 128460 301596 128512
rect 301648 128500 301654 128512
rect 306742 128500 306748 128512
rect 301648 128472 306748 128500
rect 301648 128460 301654 128472
rect 306742 128460 306748 128472
rect 306800 128460 306806 128512
rect 296070 128392 296076 128444
rect 296128 128432 296134 128444
rect 307662 128432 307668 128444
rect 296128 128404 307668 128432
rect 296128 128392 296134 128404
rect 307662 128392 307668 128404
rect 307720 128392 307726 128444
rect 178770 128324 178776 128376
rect 178828 128364 178834 128376
rect 213914 128364 213920 128376
rect 178828 128336 213920 128364
rect 178828 128324 178834 128336
rect 213914 128324 213920 128336
rect 213972 128324 213978 128376
rect 276658 128324 276664 128376
rect 276716 128364 276722 128376
rect 307570 128364 307576 128376
rect 276716 128336 307576 128364
rect 276716 128324 276722 128336
rect 307570 128324 307576 128336
rect 307628 128324 307634 128376
rect 252370 128256 252376 128308
rect 252428 128296 252434 128308
rect 282270 128296 282276 128308
rect 252428 128268 282276 128296
rect 252428 128256 252434 128268
rect 282270 128256 282276 128268
rect 282328 128256 282334 128308
rect 324314 128256 324320 128308
rect 324372 128296 324378 128308
rect 328546 128296 328552 128308
rect 324372 128268 328552 128296
rect 324372 128256 324378 128268
rect 328546 128256 328552 128268
rect 328604 128256 328610 128308
rect 252462 128188 252468 128240
rect 252520 128228 252526 128240
rect 271322 128228 271328 128240
rect 252520 128200 271328 128228
rect 252520 128188 252526 128200
rect 271322 128188 271328 128200
rect 271380 128188 271386 128240
rect 252462 127440 252468 127492
rect 252520 127480 252526 127492
rect 258902 127480 258908 127492
rect 252520 127452 258908 127480
rect 252520 127440 252526 127452
rect 258902 127440 258908 127452
rect 258960 127440 258966 127492
rect 289170 127100 289176 127152
rect 289228 127140 289234 127152
rect 307662 127140 307668 127152
rect 289228 127112 307668 127140
rect 289228 127100 289234 127112
rect 307662 127100 307668 127112
rect 307720 127100 307726 127152
rect 272518 127032 272524 127084
rect 272576 127072 272582 127084
rect 307570 127072 307576 127084
rect 272576 127044 307576 127072
rect 272576 127032 272582 127044
rect 307570 127032 307576 127044
rect 307628 127032 307634 127084
rect 271230 126964 271236 127016
rect 271288 127004 271294 127016
rect 307478 127004 307484 127016
rect 271288 126976 307484 127004
rect 271288 126964 271294 126976
rect 307478 126964 307484 126976
rect 307536 126964 307542 127016
rect 252462 126896 252468 126948
rect 252520 126936 252526 126948
rect 272610 126936 272616 126948
rect 252520 126908 272616 126936
rect 252520 126896 252526 126908
rect 272610 126896 272616 126908
rect 272668 126896 272674 126948
rect 324314 126896 324320 126948
rect 324372 126936 324378 126948
rect 328454 126936 328460 126948
rect 324372 126908 328460 126936
rect 324372 126896 324378 126908
rect 328454 126896 328460 126908
rect 328512 126896 328518 126948
rect 392578 126896 392584 126948
rect 392636 126936 392642 126948
rect 580166 126936 580172 126948
rect 392636 126908 580172 126936
rect 392636 126896 392642 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 252370 126624 252376 126676
rect 252428 126664 252434 126676
rect 258810 126664 258816 126676
rect 252428 126636 258816 126664
rect 252428 126624 252434 126636
rect 258810 126624 258816 126636
rect 258868 126624 258874 126676
rect 252186 126216 252192 126268
rect 252244 126256 252250 126268
rect 300394 126256 300400 126268
rect 252244 126228 300400 126256
rect 252244 126216 252250 126228
rect 300394 126216 300400 126228
rect 300452 126216 300458 126268
rect 300118 125740 300124 125792
rect 300176 125780 300182 125792
rect 307662 125780 307668 125792
rect 300176 125752 307668 125780
rect 300176 125740 300182 125752
rect 307662 125740 307668 125752
rect 307720 125740 307726 125792
rect 191190 125672 191196 125724
rect 191248 125712 191254 125724
rect 214006 125712 214012 125724
rect 191248 125684 214012 125712
rect 191248 125672 191254 125684
rect 214006 125672 214012 125684
rect 214064 125672 214070 125724
rect 286502 125672 286508 125724
rect 286560 125712 286566 125724
rect 307570 125712 307576 125724
rect 286560 125684 307576 125712
rect 286560 125672 286566 125684
rect 307570 125672 307576 125684
rect 307628 125672 307634 125724
rect 62022 125604 62028 125656
rect 62080 125644 62086 125656
rect 65150 125644 65156 125656
rect 62080 125616 65156 125644
rect 62080 125604 62086 125616
rect 65150 125604 65156 125616
rect 65208 125604 65214 125656
rect 169110 125604 169116 125656
rect 169168 125644 169174 125656
rect 213914 125644 213920 125656
rect 169168 125616 213920 125644
rect 169168 125604 169174 125616
rect 213914 125604 213920 125616
rect 213972 125604 213978 125656
rect 273898 125604 273904 125656
rect 273956 125644 273962 125656
rect 307478 125644 307484 125656
rect 273956 125616 307484 125644
rect 273956 125604 273962 125616
rect 307478 125604 307484 125616
rect 307536 125604 307542 125656
rect 252462 125536 252468 125588
rect 252520 125576 252526 125588
rect 274082 125576 274088 125588
rect 252520 125548 274088 125576
rect 252520 125536 252526 125548
rect 274082 125536 274088 125548
rect 274140 125536 274146 125588
rect 252370 125468 252376 125520
rect 252428 125508 252434 125520
rect 253474 125508 253480 125520
rect 252428 125480 253480 125508
rect 252428 125468 252434 125480
rect 253474 125468 253480 125480
rect 253532 125468 253538 125520
rect 275370 124924 275376 124976
rect 275428 124964 275434 124976
rect 307294 124964 307300 124976
rect 275428 124936 307300 124964
rect 275428 124924 275434 124936
rect 307294 124924 307300 124936
rect 307352 124924 307358 124976
rect 252278 124856 252284 124908
rect 252336 124896 252342 124908
rect 297450 124896 297456 124908
rect 252336 124868 297456 124896
rect 252336 124856 252342 124868
rect 297450 124856 297456 124868
rect 297508 124856 297514 124908
rect 303062 124312 303068 124364
rect 303120 124352 303126 124364
rect 306926 124352 306932 124364
rect 303120 124324 306932 124352
rect 303120 124312 303126 124324
rect 306926 124312 306932 124324
rect 306984 124312 306990 124364
rect 180058 124244 180064 124296
rect 180116 124284 180122 124296
rect 213914 124284 213920 124296
rect 180116 124256 213920 124284
rect 180116 124244 180122 124256
rect 213914 124244 213920 124256
rect 213972 124244 213978 124296
rect 298922 124244 298928 124296
rect 298980 124284 298986 124296
rect 307570 124284 307576 124296
rect 298980 124256 307576 124284
rect 298980 124244 298986 124256
rect 307570 124244 307576 124256
rect 307628 124244 307634 124296
rect 170582 124176 170588 124228
rect 170640 124216 170646 124228
rect 214006 124216 214012 124228
rect 170640 124188 214012 124216
rect 170640 124176 170646 124188
rect 214006 124176 214012 124188
rect 214064 124176 214070 124228
rect 295978 124176 295984 124228
rect 296036 124216 296042 124228
rect 307662 124216 307668 124228
rect 296036 124188 307668 124216
rect 296036 124176 296042 124188
rect 307662 124176 307668 124188
rect 307720 124176 307726 124228
rect 252462 124108 252468 124160
rect 252520 124148 252526 124160
rect 269758 124148 269764 124160
rect 252520 124120 269764 124148
rect 252520 124108 252526 124120
rect 269758 124108 269764 124120
rect 269816 124108 269822 124160
rect 324314 124108 324320 124160
rect 324372 124148 324378 124160
rect 340874 124148 340880 124160
rect 324372 124120 340880 124148
rect 324372 124108 324378 124120
rect 340874 124108 340880 124120
rect 340932 124108 340938 124160
rect 252370 124040 252376 124092
rect 252428 124080 252434 124092
rect 261478 124080 261484 124092
rect 252428 124052 261484 124080
rect 252428 124040 252434 124052
rect 261478 124040 261484 124052
rect 261536 124040 261542 124092
rect 252278 123428 252284 123480
rect 252336 123468 252342 123480
rect 304534 123468 304540 123480
rect 252336 123440 304540 123468
rect 252336 123428 252342 123440
rect 304534 123428 304540 123440
rect 304592 123428 304598 123480
rect 211798 123360 211804 123412
rect 211856 123400 211862 123412
rect 213914 123400 213920 123412
rect 211856 123372 213920 123400
rect 211856 123360 211862 123372
rect 213914 123360 213920 123372
rect 213972 123360 213978 123412
rect 304350 122952 304356 123004
rect 304408 122992 304414 123004
rect 307662 122992 307668 123004
rect 304408 122964 307668 122992
rect 304408 122952 304414 122964
rect 307662 122952 307668 122964
rect 307720 122952 307726 123004
rect 292022 122884 292028 122936
rect 292080 122924 292086 122936
rect 307478 122924 307484 122936
rect 292080 122896 307484 122924
rect 292080 122884 292086 122896
rect 307478 122884 307484 122896
rect 307536 122884 307542 122936
rect 195330 122816 195336 122868
rect 195388 122856 195394 122868
rect 213914 122856 213920 122868
rect 195388 122828 213920 122856
rect 195388 122816 195394 122828
rect 213914 122816 213920 122828
rect 213972 122816 213978 122868
rect 282362 122816 282368 122868
rect 282420 122856 282426 122868
rect 307570 122856 307576 122868
rect 282420 122828 307576 122856
rect 282420 122816 282426 122828
rect 307570 122816 307576 122828
rect 307628 122816 307634 122868
rect 324314 122748 324320 122800
rect 324372 122788 324378 122800
rect 336734 122788 336740 122800
rect 324372 122760 336740 122788
rect 324372 122748 324378 122760
rect 336734 122748 336740 122760
rect 336792 122748 336798 122800
rect 252370 122680 252376 122732
rect 252428 122720 252434 122732
rect 286318 122720 286324 122732
rect 252428 122692 286324 122720
rect 252428 122680 252434 122692
rect 286318 122680 286324 122692
rect 286376 122680 286382 122732
rect 252462 122612 252468 122664
rect 252520 122652 252526 122664
rect 289354 122652 289360 122664
rect 252520 122624 289360 122652
rect 252520 122612 252526 122624
rect 289354 122612 289360 122624
rect 289412 122612 289418 122664
rect 297542 121592 297548 121644
rect 297600 121632 297606 121644
rect 307570 121632 307576 121644
rect 297600 121604 307576 121632
rect 297600 121592 297606 121604
rect 307570 121592 307576 121604
rect 307628 121592 307634 121644
rect 202230 121524 202236 121576
rect 202288 121564 202294 121576
rect 213914 121564 213920 121576
rect 202288 121536 213920 121564
rect 202288 121524 202294 121536
rect 213914 121524 213920 121536
rect 213972 121524 213978 121576
rect 289262 121524 289268 121576
rect 289320 121564 289326 121576
rect 307662 121564 307668 121576
rect 289320 121536 307668 121564
rect 289320 121524 289326 121536
rect 307662 121524 307668 121536
rect 307720 121524 307726 121576
rect 182818 121456 182824 121508
rect 182876 121496 182882 121508
rect 214006 121496 214012 121508
rect 182876 121468 214012 121496
rect 182876 121456 182882 121468
rect 214006 121456 214012 121468
rect 214064 121456 214070 121508
rect 286410 121456 286416 121508
rect 286468 121496 286474 121508
rect 307478 121496 307484 121508
rect 286468 121468 307484 121496
rect 286468 121456 286474 121468
rect 307478 121456 307484 121468
rect 307536 121456 307542 121508
rect 252370 121388 252376 121440
rect 252428 121428 252434 121440
rect 290642 121428 290648 121440
rect 252428 121400 290648 121428
rect 252428 121388 252434 121400
rect 290642 121388 290648 121400
rect 290700 121388 290706 121440
rect 324406 121388 324412 121440
rect 324464 121428 324470 121440
rect 343818 121428 343824 121440
rect 324464 121400 343824 121428
rect 324464 121388 324470 121400
rect 343818 121388 343824 121400
rect 343876 121388 343882 121440
rect 324314 121320 324320 121372
rect 324372 121360 324378 121372
rect 338298 121360 338304 121372
rect 324372 121332 338304 121360
rect 324372 121320 324378 121332
rect 338298 121320 338304 121332
rect 338356 121320 338362 121372
rect 251910 120708 251916 120760
rect 251968 120748 251974 120760
rect 268470 120748 268476 120760
rect 251968 120720 268476 120748
rect 251968 120708 251974 120720
rect 268470 120708 268476 120720
rect 268528 120708 268534 120760
rect 252462 120640 252468 120692
rect 252520 120680 252526 120692
rect 260098 120680 260104 120692
rect 252520 120652 260104 120680
rect 252520 120640 252526 120652
rect 260098 120640 260104 120652
rect 260156 120640 260162 120692
rect 291838 120232 291844 120284
rect 291896 120272 291902 120284
rect 307662 120272 307668 120284
rect 291896 120244 307668 120272
rect 291896 120232 291902 120244
rect 307662 120232 307668 120244
rect 307720 120232 307726 120284
rect 290458 120164 290464 120216
rect 290516 120204 290522 120216
rect 307570 120204 307576 120216
rect 290516 120176 307576 120204
rect 290516 120164 290522 120176
rect 307570 120164 307576 120176
rect 307628 120164 307634 120216
rect 170674 120096 170680 120148
rect 170732 120136 170738 120148
rect 213914 120136 213920 120148
rect 170732 120108 213920 120136
rect 170732 120096 170738 120108
rect 213914 120096 213920 120108
rect 213972 120096 213978 120148
rect 269758 120096 269764 120148
rect 269816 120136 269822 120148
rect 307478 120136 307484 120148
rect 269816 120108 307484 120136
rect 269816 120096 269822 120108
rect 307478 120096 307484 120108
rect 307536 120096 307542 120148
rect 252370 120028 252376 120080
rect 252428 120068 252434 120080
rect 298738 120068 298744 120080
rect 252428 120040 298744 120068
rect 252428 120028 252434 120040
rect 298738 120028 298744 120040
rect 298796 120028 298802 120080
rect 324314 120028 324320 120080
rect 324372 120068 324378 120080
rect 338206 120068 338212 120080
rect 324372 120040 338212 120068
rect 324372 120028 324378 120040
rect 338206 120028 338212 120040
rect 338264 120028 338270 120080
rect 252462 119960 252468 120012
rect 252520 120000 252526 120012
rect 262950 120000 262956 120012
rect 252520 119972 262956 120000
rect 252520 119960 252526 119972
rect 262950 119960 262956 119972
rect 263008 119960 263014 120012
rect 252462 119416 252468 119468
rect 252520 119456 252526 119468
rect 258718 119456 258724 119468
rect 252520 119428 258724 119456
rect 252520 119416 252526 119428
rect 258718 119416 258724 119428
rect 258776 119416 258782 119468
rect 263042 119348 263048 119400
rect 263100 119388 263106 119400
rect 307386 119388 307392 119400
rect 263100 119360 307392 119388
rect 263100 119348 263106 119360
rect 307386 119348 307392 119360
rect 307444 119348 307450 119400
rect 178862 118804 178868 118856
rect 178920 118844 178926 118856
rect 214006 118844 214012 118856
rect 178920 118816 214012 118844
rect 178920 118804 178926 118816
rect 214006 118804 214012 118816
rect 214064 118804 214070 118856
rect 298830 118804 298836 118856
rect 298888 118844 298894 118856
rect 307662 118844 307668 118856
rect 298888 118816 307668 118844
rect 298888 118804 298894 118816
rect 307662 118804 307668 118816
rect 307720 118804 307726 118856
rect 172054 118736 172060 118788
rect 172112 118776 172118 118788
rect 214098 118776 214104 118788
rect 172112 118748 214104 118776
rect 172112 118736 172118 118748
rect 214098 118736 214104 118748
rect 214156 118736 214162 118788
rect 167914 118668 167920 118720
rect 167972 118708 167978 118720
rect 213914 118708 213920 118720
rect 167972 118680 213920 118708
rect 167972 118668 167978 118680
rect 213914 118668 213920 118680
rect 213972 118668 213978 118720
rect 301682 118668 301688 118720
rect 301740 118708 301746 118720
rect 307478 118708 307484 118720
rect 301740 118680 307484 118708
rect 301740 118668 301746 118680
rect 307478 118668 307484 118680
rect 307536 118668 307542 118720
rect 252462 118600 252468 118652
rect 252520 118640 252526 118652
rect 267090 118640 267096 118652
rect 252520 118612 267096 118640
rect 252520 118600 252526 118612
rect 267090 118600 267096 118612
rect 267148 118600 267154 118652
rect 324314 118600 324320 118652
rect 324372 118640 324378 118652
rect 340966 118640 340972 118652
rect 324372 118612 340972 118640
rect 324372 118600 324378 118612
rect 340966 118600 340972 118612
rect 341024 118600 341030 118652
rect 252370 118532 252376 118584
rect 252428 118572 252434 118584
rect 256142 118572 256148 118584
rect 252428 118544 256148 118572
rect 252428 118532 252434 118544
rect 256142 118532 256148 118544
rect 256200 118532 256206 118584
rect 324406 118532 324412 118584
rect 324464 118572 324470 118584
rect 332686 118572 332692 118584
rect 324464 118544 332692 118572
rect 324464 118532 324470 118544
rect 332686 118532 332692 118544
rect 332744 118532 332750 118584
rect 174722 117920 174728 117972
rect 174780 117960 174786 117972
rect 214742 117960 214748 117972
rect 174780 117932 214748 117960
rect 174780 117920 174786 117932
rect 214742 117920 214748 117932
rect 214800 117920 214806 117972
rect 252278 117920 252284 117972
rect 252336 117960 252342 117972
rect 296162 117960 296168 117972
rect 252336 117932 296168 117960
rect 252336 117920 252342 117932
rect 296162 117920 296168 117932
rect 296220 117920 296226 117972
rect 293310 117444 293316 117496
rect 293368 117484 293374 117496
rect 307662 117484 307668 117496
rect 293368 117456 307668 117484
rect 293368 117444 293374 117456
rect 307662 117444 307668 117456
rect 307720 117444 307726 117496
rect 268378 117376 268384 117428
rect 268436 117416 268442 117428
rect 307570 117416 307576 117428
rect 268436 117388 307576 117416
rect 268436 117376 268442 117388
rect 307570 117376 307576 117388
rect 307628 117376 307634 117428
rect 181438 117308 181444 117360
rect 181496 117348 181502 117360
rect 213914 117348 213920 117360
rect 181496 117320 213920 117348
rect 181496 117308 181502 117320
rect 213914 117308 213920 117320
rect 213972 117308 213978 117360
rect 260098 117308 260104 117360
rect 260156 117348 260162 117360
rect 306558 117348 306564 117360
rect 260156 117320 306564 117348
rect 260156 117308 260162 117320
rect 306558 117308 306564 117320
rect 306616 117308 306622 117360
rect 252462 117240 252468 117292
rect 252520 117280 252526 117292
rect 262858 117280 262864 117292
rect 252520 117252 262864 117280
rect 252520 117240 252526 117252
rect 262858 117240 262864 117252
rect 262916 117240 262922 117292
rect 324314 117240 324320 117292
rect 324372 117280 324378 117292
rect 333974 117280 333980 117292
rect 324372 117252 333980 117280
rect 324372 117240 324378 117252
rect 333974 117240 333980 117252
rect 334032 117240 334038 117292
rect 252094 116560 252100 116612
rect 252152 116600 252158 116612
rect 281074 116600 281080 116612
rect 252152 116572 281080 116600
rect 252152 116560 252158 116572
rect 281074 116560 281080 116572
rect 281132 116560 281138 116612
rect 252462 116084 252468 116136
rect 252520 116124 252526 116136
rect 260190 116124 260196 116136
rect 252520 116096 260196 116124
rect 252520 116084 252526 116096
rect 260190 116084 260196 116096
rect 260248 116084 260254 116136
rect 296162 116084 296168 116136
rect 296220 116124 296226 116136
rect 307570 116124 307576 116136
rect 296220 116096 307576 116124
rect 296220 116084 296226 116096
rect 307570 116084 307576 116096
rect 307628 116084 307634 116136
rect 186958 116016 186964 116068
rect 187016 116056 187022 116068
rect 213914 116056 213920 116068
rect 187016 116028 213920 116056
rect 187016 116016 187022 116028
rect 213914 116016 213920 116028
rect 213972 116016 213978 116068
rect 280890 116016 280896 116068
rect 280948 116056 280954 116068
rect 307662 116056 307668 116068
rect 280948 116028 307668 116056
rect 280948 116016 280954 116028
rect 307662 116016 307668 116028
rect 307720 116016 307726 116068
rect 176102 115948 176108 116000
rect 176160 115988 176166 116000
rect 214006 115988 214012 116000
rect 176160 115960 214012 115988
rect 176160 115948 176166 115960
rect 214006 115948 214012 115960
rect 214064 115948 214070 116000
rect 267182 115948 267188 116000
rect 267240 115988 267246 116000
rect 306742 115988 306748 116000
rect 267240 115960 306748 115988
rect 267240 115948 267246 115960
rect 306742 115948 306748 115960
rect 306800 115948 306806 116000
rect 252370 115880 252376 115932
rect 252428 115920 252434 115932
rect 264514 115920 264520 115932
rect 252428 115892 264520 115920
rect 252428 115880 252434 115892
rect 264514 115880 264520 115892
rect 264572 115880 264578 115932
rect 252278 115200 252284 115252
rect 252336 115240 252342 115252
rect 282454 115240 282460 115252
rect 252336 115212 282460 115240
rect 252336 115200 252342 115212
rect 282454 115200 282460 115212
rect 282512 115200 282518 115252
rect 293402 114656 293408 114708
rect 293460 114696 293466 114708
rect 307570 114696 307576 114708
rect 293460 114668 307576 114696
rect 293460 114656 293466 114668
rect 307570 114656 307576 114668
rect 307628 114656 307634 114708
rect 180150 114588 180156 114640
rect 180208 114628 180214 114640
rect 213914 114628 213920 114640
rect 180208 114600 213920 114628
rect 180208 114588 180214 114600
rect 213914 114588 213920 114600
rect 213972 114588 213978 114640
rect 287882 114588 287888 114640
rect 287940 114628 287946 114640
rect 307662 114628 307668 114640
rect 287940 114600 307668 114628
rect 287940 114588 287946 114600
rect 307662 114588 307668 114600
rect 307720 114588 307726 114640
rect 176010 114520 176016 114572
rect 176068 114560 176074 114572
rect 214006 114560 214012 114572
rect 176068 114532 214012 114560
rect 176068 114520 176074 114532
rect 214006 114520 214012 114532
rect 214064 114520 214070 114572
rect 264238 114520 264244 114572
rect 264296 114560 264302 114572
rect 307478 114560 307484 114572
rect 264296 114532 307484 114560
rect 264296 114520 264302 114532
rect 307478 114520 307484 114532
rect 307536 114520 307542 114572
rect 252462 114452 252468 114504
rect 252520 114492 252526 114504
rect 300210 114492 300216 114504
rect 252520 114464 300216 114492
rect 252520 114452 252526 114464
rect 300210 114452 300216 114464
rect 300268 114452 300274 114504
rect 324314 114452 324320 114504
rect 324372 114492 324378 114504
rect 342346 114492 342352 114504
rect 324372 114464 342352 114492
rect 324372 114452 324378 114464
rect 342346 114452 342352 114464
rect 342404 114452 342410 114504
rect 252370 114384 252376 114436
rect 252428 114424 252434 114436
rect 285030 114424 285036 114436
rect 252428 114396 285036 114424
rect 252428 114384 252434 114396
rect 285030 114384 285036 114396
rect 285088 114384 285094 114436
rect 324406 114384 324412 114436
rect 324464 114424 324470 114436
rect 335538 114424 335544 114436
rect 324464 114396 335544 114424
rect 324464 114384 324470 114396
rect 335538 114384 335544 114396
rect 335596 114384 335602 114436
rect 211890 113228 211896 113280
rect 211948 113268 211954 113280
rect 214006 113268 214012 113280
rect 211948 113240 214012 113268
rect 211948 113228 211954 113240
rect 214006 113228 214012 113240
rect 214064 113228 214070 113280
rect 294598 113228 294604 113280
rect 294656 113268 294662 113280
rect 307662 113268 307668 113280
rect 294656 113240 307668 113268
rect 294656 113228 294662 113240
rect 307662 113228 307668 113240
rect 307720 113228 307726 113280
rect 198090 113160 198096 113212
rect 198148 113200 198154 113212
rect 213914 113200 213920 113212
rect 198148 113172 213920 113200
rect 198148 113160 198154 113172
rect 213914 113160 213920 113172
rect 213972 113160 213978 113212
rect 284938 113160 284944 113212
rect 284996 113200 285002 113212
rect 307570 113200 307576 113212
rect 284996 113172 307576 113200
rect 284996 113160 285002 113172
rect 307570 113160 307576 113172
rect 307628 113160 307634 113212
rect 252462 113092 252468 113144
rect 252520 113132 252526 113144
rect 299106 113132 299112 113144
rect 252520 113104 299112 113132
rect 252520 113092 252526 113104
rect 299106 113092 299112 113104
rect 299164 113092 299170 113144
rect 324314 113092 324320 113144
rect 324372 113132 324378 113144
rect 337010 113132 337016 113144
rect 324372 113104 337016 113132
rect 324372 113092 324378 113104
rect 337010 113092 337016 113104
rect 337068 113092 337074 113144
rect 252002 112412 252008 112464
rect 252060 112452 252066 112464
rect 305638 112452 305644 112464
rect 252060 112424 305644 112452
rect 252060 112412 252066 112424
rect 305638 112412 305644 112424
rect 305696 112412 305702 112464
rect 204990 111868 204996 111920
rect 205048 111908 205054 111920
rect 214006 111908 214012 111920
rect 205048 111880 214012 111908
rect 205048 111868 205054 111880
rect 214006 111868 214012 111880
rect 214064 111868 214070 111920
rect 301498 111868 301504 111920
rect 301556 111908 301562 111920
rect 307478 111908 307484 111920
rect 301556 111880 307484 111908
rect 301556 111868 301562 111880
rect 307478 111868 307484 111880
rect 307536 111868 307542 111920
rect 169202 111800 169208 111852
rect 169260 111840 169266 111852
rect 213914 111840 213920 111852
rect 169260 111812 213920 111840
rect 169260 111800 169266 111812
rect 213914 111800 213920 111812
rect 213972 111800 213978 111852
rect 253198 111800 253204 111852
rect 253256 111840 253262 111852
rect 307662 111840 307668 111852
rect 253256 111812 307668 111840
rect 253256 111800 253262 111812
rect 307662 111800 307668 111812
rect 307720 111800 307726 111852
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 17218 111772 17224 111784
rect 3200 111744 17224 111772
rect 3200 111732 3206 111744
rect 17218 111732 17224 111744
rect 17276 111732 17282 111784
rect 168006 111732 168012 111784
rect 168064 111772 168070 111784
rect 171962 111772 171968 111784
rect 168064 111744 171968 111772
rect 168064 111732 168070 111744
rect 171962 111732 171968 111744
rect 172020 111732 172026 111784
rect 252462 111732 252468 111784
rect 252520 111772 252526 111784
rect 304258 111772 304264 111784
rect 252520 111744 304264 111772
rect 252520 111732 252526 111744
rect 304258 111732 304264 111744
rect 304316 111732 304322 111784
rect 252370 111664 252376 111716
rect 252428 111704 252434 111716
rect 256050 111704 256056 111716
rect 252428 111676 256056 111704
rect 252428 111664 252434 111676
rect 256050 111664 256056 111676
rect 256108 111664 256114 111716
rect 252278 111052 252284 111104
rect 252336 111092 252342 111104
rect 301774 111092 301780 111104
rect 252336 111064 301780 111092
rect 252336 111052 252342 111064
rect 301774 111052 301780 111064
rect 301832 111052 301838 111104
rect 192478 110508 192484 110560
rect 192536 110548 192542 110560
rect 214006 110548 214012 110560
rect 192536 110520 214012 110548
rect 192536 110508 192542 110520
rect 214006 110508 214012 110520
rect 214064 110508 214070 110560
rect 300210 110508 300216 110560
rect 300268 110548 300274 110560
rect 307570 110548 307576 110560
rect 300268 110520 307576 110548
rect 300268 110508 300274 110520
rect 307570 110508 307576 110520
rect 307628 110508 307634 110560
rect 173434 110440 173440 110492
rect 173492 110480 173498 110492
rect 213914 110480 213920 110492
rect 173492 110452 213920 110480
rect 173492 110440 173498 110452
rect 213914 110440 213920 110452
rect 213972 110440 213978 110492
rect 303154 110440 303160 110492
rect 303212 110480 303218 110492
rect 307662 110480 307668 110492
rect 303212 110452 307668 110480
rect 303212 110440 303218 110452
rect 307662 110440 307668 110452
rect 307720 110440 307726 110492
rect 168098 110372 168104 110424
rect 168156 110412 168162 110424
rect 175918 110412 175924 110424
rect 168156 110384 175924 110412
rect 168156 110372 168162 110384
rect 175918 110372 175924 110384
rect 175976 110372 175982 110424
rect 252370 110372 252376 110424
rect 252428 110412 252434 110424
rect 287974 110412 287980 110424
rect 252428 110384 287980 110412
rect 252428 110372 252434 110384
rect 287974 110372 287980 110384
rect 288032 110372 288038 110424
rect 252462 110304 252468 110356
rect 252520 110344 252526 110356
rect 264330 110344 264336 110356
rect 252520 110316 264336 110344
rect 252520 110304 252526 110316
rect 264330 110304 264336 110316
rect 264388 110304 264394 110356
rect 251634 110236 251640 110288
rect 251692 110276 251698 110288
rect 254578 110276 254584 110288
rect 251692 110248 254584 110276
rect 251692 110236 251698 110248
rect 254578 110236 254584 110248
rect 254636 110236 254642 110288
rect 304534 109148 304540 109200
rect 304592 109188 304598 109200
rect 307478 109188 307484 109200
rect 304592 109160 307484 109188
rect 304592 109148 304598 109160
rect 307478 109148 307484 109160
rect 307536 109148 307542 109200
rect 209130 109080 209136 109132
rect 209188 109120 209194 109132
rect 214006 109120 214012 109132
rect 209188 109092 214012 109120
rect 209188 109080 209194 109092
rect 214006 109080 214012 109092
rect 214064 109080 214070 109132
rect 287790 109080 287796 109132
rect 287848 109120 287854 109132
rect 307570 109120 307576 109132
rect 287848 109092 307576 109120
rect 287848 109080 287854 109092
rect 307570 109080 307576 109092
rect 307628 109080 307634 109132
rect 174630 109012 174636 109064
rect 174688 109052 174694 109064
rect 213914 109052 213920 109064
rect 174688 109024 213920 109052
rect 174688 109012 174694 109024
rect 213914 109012 213920 109024
rect 213972 109012 213978 109064
rect 262858 109012 262864 109064
rect 262916 109052 262922 109064
rect 307662 109052 307668 109064
rect 262916 109024 307668 109052
rect 262916 109012 262922 109024
rect 307662 109012 307668 109024
rect 307720 109012 307726 109064
rect 168006 108944 168012 108996
rect 168064 108984 168070 108996
rect 177574 108984 177580 108996
rect 168064 108956 177580 108984
rect 168064 108944 168070 108956
rect 177574 108944 177580 108956
rect 177632 108944 177638 108996
rect 252370 108944 252376 108996
rect 252428 108984 252434 108996
rect 292114 108984 292120 108996
rect 252428 108956 292120 108984
rect 252428 108944 252434 108956
rect 292114 108944 292120 108956
rect 292172 108944 292178 108996
rect 324314 108944 324320 108996
rect 324372 108984 324378 108996
rect 353294 108984 353300 108996
rect 324372 108956 353300 108984
rect 324372 108944 324378 108956
rect 353294 108944 353300 108956
rect 353352 108944 353358 108996
rect 252462 108876 252468 108928
rect 252520 108916 252526 108928
rect 275370 108916 275376 108928
rect 252520 108888 275376 108916
rect 252520 108876 252526 108888
rect 275370 108876 275376 108888
rect 275428 108876 275434 108928
rect 282270 107856 282276 107908
rect 282328 107896 282334 107908
rect 307662 107896 307668 107908
rect 282328 107868 307668 107896
rect 282328 107856 282334 107868
rect 307662 107856 307668 107868
rect 307720 107856 307726 107908
rect 292206 107720 292212 107772
rect 292264 107760 292270 107772
rect 307662 107760 307668 107772
rect 292264 107732 307668 107760
rect 292264 107720 292270 107732
rect 307662 107720 307668 107732
rect 307720 107720 307726 107772
rect 177666 107652 177672 107704
rect 177724 107692 177730 107704
rect 213914 107692 213920 107704
rect 177724 107664 213920 107692
rect 177724 107652 177730 107664
rect 213914 107652 213920 107664
rect 213972 107652 213978 107704
rect 302970 107652 302976 107704
rect 303028 107692 303034 107704
rect 307570 107692 307576 107704
rect 303028 107664 307576 107692
rect 303028 107652 303034 107664
rect 307570 107652 307576 107664
rect 307628 107652 307634 107704
rect 252370 107584 252376 107636
rect 252428 107624 252434 107636
rect 305914 107624 305920 107636
rect 252428 107596 305920 107624
rect 252428 107584 252434 107596
rect 305914 107584 305920 107596
rect 305972 107584 305978 107636
rect 252462 107516 252468 107568
rect 252520 107556 252526 107568
rect 264422 107556 264428 107568
rect 252520 107528 264428 107556
rect 252520 107516 252526 107528
rect 264422 107516 264428 107528
rect 264480 107516 264486 107568
rect 252186 107448 252192 107500
rect 252244 107488 252250 107500
rect 254670 107488 254676 107500
rect 252244 107460 254676 107488
rect 252244 107448 252250 107460
rect 254670 107448 254676 107460
rect 254728 107448 254734 107500
rect 268470 106428 268476 106480
rect 268528 106468 268534 106480
rect 307478 106468 307484 106480
rect 268528 106440 307484 106468
rect 268528 106428 268534 106440
rect 307478 106428 307484 106440
rect 307536 106428 307542 106480
rect 304258 106360 304264 106412
rect 304316 106400 304322 106412
rect 307662 106400 307668 106412
rect 304316 106372 307668 106400
rect 304316 106360 304322 106372
rect 307662 106360 307668 106372
rect 307720 106360 307726 106412
rect 169294 106292 169300 106344
rect 169352 106332 169358 106344
rect 213914 106332 213920 106344
rect 169352 106304 213920 106332
rect 169352 106292 169358 106304
rect 213914 106292 213920 106304
rect 213972 106292 213978 106344
rect 252462 106224 252468 106276
rect 252520 106264 252526 106276
rect 285214 106264 285220 106276
rect 252520 106236 285220 106264
rect 252520 106224 252526 106236
rect 285214 106224 285220 106236
rect 285272 106224 285278 106276
rect 252278 106156 252284 106208
rect 252336 106196 252342 106208
rect 255958 106196 255964 106208
rect 252336 106168 255964 106196
rect 252336 106156 252342 106168
rect 255958 106156 255964 106168
rect 256016 106156 256022 106208
rect 252370 105544 252376 105596
rect 252428 105584 252434 105596
rect 299014 105584 299020 105596
rect 252428 105556 299020 105584
rect 252428 105544 252434 105556
rect 299014 105544 299020 105556
rect 299072 105544 299078 105596
rect 300486 105000 300492 105052
rect 300544 105040 300550 105052
rect 307662 105040 307668 105052
rect 300544 105012 307668 105040
rect 300544 105000 300550 105012
rect 307662 105000 307668 105012
rect 307720 105000 307726 105052
rect 207750 104932 207756 104984
rect 207808 104972 207814 104984
rect 213914 104972 213920 104984
rect 207808 104944 213920 104972
rect 207808 104932 207814 104944
rect 213914 104932 213920 104944
rect 213972 104932 213978 104984
rect 298738 104932 298744 104984
rect 298796 104972 298802 104984
rect 307478 104972 307484 104984
rect 298796 104944 307484 104972
rect 298796 104932 298802 104944
rect 307478 104932 307484 104944
rect 307536 104932 307542 104984
rect 199470 104864 199476 104916
rect 199528 104904 199534 104916
rect 214006 104904 214012 104916
rect 199528 104876 214012 104904
rect 199528 104864 199534 104876
rect 214006 104864 214012 104876
rect 214064 104864 214070 104916
rect 285030 104864 285036 104916
rect 285088 104904 285094 104916
rect 307570 104904 307576 104916
rect 285088 104876 307576 104904
rect 285088 104864 285094 104876
rect 307570 104864 307576 104876
rect 307628 104864 307634 104916
rect 252462 104796 252468 104848
rect 252520 104836 252526 104848
rect 265618 104836 265624 104848
rect 252520 104808 265624 104836
rect 252520 104796 252526 104808
rect 265618 104796 265624 104808
rect 265676 104796 265682 104848
rect 252278 104728 252284 104780
rect 252336 104768 252342 104780
rect 257430 104768 257436 104780
rect 252336 104740 257436 104768
rect 252336 104728 252342 104740
rect 257430 104728 257436 104740
rect 257488 104728 257494 104780
rect 251266 104116 251272 104168
rect 251324 104156 251330 104168
rect 275278 104156 275284 104168
rect 251324 104128 275284 104156
rect 251324 104116 251330 104128
rect 275278 104116 275284 104128
rect 275336 104116 275342 104168
rect 210602 103844 210608 103896
rect 210660 103884 210666 103896
rect 213914 103884 213920 103896
rect 210660 103856 213920 103884
rect 210660 103844 210666 103856
rect 213914 103844 213920 103856
rect 213972 103844 213978 103896
rect 279418 103572 279424 103624
rect 279476 103612 279482 103624
rect 307662 103612 307668 103624
rect 279476 103584 307668 103612
rect 279476 103572 279482 103584
rect 307662 103572 307668 103584
rect 307720 103572 307726 103624
rect 171962 103504 171968 103556
rect 172020 103544 172026 103556
rect 213914 103544 213920 103556
rect 172020 103516 213920 103544
rect 172020 103504 172026 103516
rect 213914 103504 213920 103516
rect 213972 103504 213978 103556
rect 267090 103504 267096 103556
rect 267148 103544 267154 103556
rect 307570 103544 307576 103556
rect 267148 103516 307576 103544
rect 267148 103504 267154 103516
rect 307570 103504 307576 103516
rect 307628 103504 307634 103556
rect 252462 103436 252468 103488
rect 252520 103476 252526 103488
rect 268562 103476 268568 103488
rect 252520 103448 268568 103476
rect 252520 103436 252526 103448
rect 268562 103436 268568 103448
rect 268620 103436 268626 103488
rect 324406 103436 324412 103488
rect 324464 103476 324470 103488
rect 339678 103476 339684 103488
rect 324464 103448 339684 103476
rect 324464 103436 324470 103448
rect 339678 103436 339684 103448
rect 339736 103436 339742 103488
rect 251174 103300 251180 103352
rect 251232 103340 251238 103352
rect 253382 103340 253388 103352
rect 251232 103312 253388 103340
rect 251232 103300 251238 103312
rect 253382 103300 253388 103312
rect 253440 103300 253446 103352
rect 252186 102756 252192 102808
rect 252244 102796 252250 102808
rect 269942 102796 269948 102808
rect 252244 102768 269948 102796
rect 252244 102756 252250 102768
rect 269942 102756 269948 102768
rect 270000 102756 270006 102808
rect 294690 102280 294696 102332
rect 294748 102320 294754 102332
rect 306926 102320 306932 102332
rect 294748 102292 306932 102320
rect 294748 102280 294754 102292
rect 306926 102280 306932 102292
rect 306984 102280 306990 102332
rect 275278 102212 275284 102264
rect 275336 102252 275342 102264
rect 307570 102252 307576 102264
rect 275336 102224 307576 102252
rect 275336 102212 275342 102224
rect 307570 102212 307576 102224
rect 307628 102212 307634 102264
rect 269850 102144 269856 102196
rect 269908 102184 269914 102196
rect 307662 102184 307668 102196
rect 269908 102156 307668 102184
rect 269908 102144 269914 102156
rect 307662 102144 307668 102156
rect 307720 102144 307726 102196
rect 251358 102076 251364 102128
rect 251416 102116 251422 102128
rect 253290 102116 253296 102128
rect 251416 102088 253296 102116
rect 251416 102076 251422 102088
rect 253290 102076 253296 102088
rect 253348 102076 253354 102128
rect 252462 102008 252468 102060
rect 252520 102048 252526 102060
rect 280982 102048 280988 102060
rect 252520 102020 280988 102048
rect 252520 102008 252526 102020
rect 280982 102008 280988 102020
rect 281040 102008 281046 102060
rect 252278 101396 252284 101448
rect 252336 101436 252342 101448
rect 300302 101436 300308 101448
rect 252336 101408 300308 101436
rect 252336 101396 252342 101408
rect 300302 101396 300308 101408
rect 300360 101396 300366 101448
rect 300394 100852 300400 100904
rect 300452 100892 300458 100904
rect 307570 100892 307576 100904
rect 300452 100864 307576 100892
rect 300452 100852 300458 100864
rect 307570 100852 307576 100864
rect 307628 100852 307634 100904
rect 299014 100784 299020 100836
rect 299072 100824 299078 100836
rect 307478 100824 307484 100836
rect 299072 100796 307484 100824
rect 299072 100784 299078 100796
rect 307478 100784 307484 100796
rect 307536 100784 307542 100836
rect 283650 100716 283656 100768
rect 283708 100756 283714 100768
rect 307662 100756 307668 100768
rect 283708 100728 307668 100756
rect 283708 100716 283714 100728
rect 307662 100716 307668 100728
rect 307720 100716 307726 100768
rect 252370 100648 252376 100700
rect 252428 100688 252434 100700
rect 304442 100688 304448 100700
rect 252428 100660 304448 100688
rect 252428 100648 252434 100660
rect 304442 100648 304448 100660
rect 304500 100648 304506 100700
rect 252462 100580 252468 100632
rect 252520 100620 252526 100632
rect 294874 100620 294880 100632
rect 252520 100592 294880 100620
rect 252520 100580 252526 100592
rect 294874 100580 294880 100592
rect 294932 100580 294938 100632
rect 166534 99424 166540 99476
rect 166592 99464 166598 99476
rect 213914 99464 213920 99476
rect 166592 99436 213920 99464
rect 166592 99424 166598 99436
rect 213914 99424 213920 99436
rect 213972 99424 213978 99476
rect 297450 99424 297456 99476
rect 297508 99464 297514 99476
rect 307570 99464 307576 99476
rect 297508 99436 307576 99464
rect 297508 99424 297514 99436
rect 307570 99424 307576 99436
rect 307628 99424 307634 99476
rect 166350 99356 166356 99408
rect 166408 99396 166414 99408
rect 214006 99396 214012 99408
rect 166408 99368 214012 99396
rect 166408 99356 166414 99368
rect 214006 99356 214012 99368
rect 214064 99356 214070 99408
rect 290642 99356 290648 99408
rect 290700 99396 290706 99408
rect 307662 99396 307668 99408
rect 290700 99368 307668 99396
rect 290700 99356 290706 99368
rect 307662 99356 307668 99368
rect 307720 99356 307726 99408
rect 252370 99288 252376 99340
rect 252428 99328 252434 99340
rect 286594 99328 286600 99340
rect 252428 99300 286600 99328
rect 252428 99288 252434 99300
rect 286594 99288 286600 99300
rect 286652 99288 286658 99340
rect 252462 99220 252468 99272
rect 252520 99260 252526 99272
rect 257338 99260 257344 99272
rect 252520 99232 257344 99260
rect 252520 99220 252526 99232
rect 257338 99220 257344 99232
rect 257396 99220 257402 99272
rect 166442 98064 166448 98116
rect 166500 98104 166506 98116
rect 214006 98104 214012 98116
rect 166500 98076 214012 98104
rect 166500 98064 166506 98076
rect 214006 98064 214012 98076
rect 214064 98064 214070 98116
rect 286318 98064 286324 98116
rect 286376 98104 286382 98116
rect 307570 98104 307576 98116
rect 286376 98076 307576 98104
rect 286376 98064 286382 98076
rect 307570 98064 307576 98076
rect 307628 98064 307634 98116
rect 164970 97996 164976 98048
rect 165028 98036 165034 98048
rect 213914 98036 213920 98048
rect 165028 98008 213920 98036
rect 165028 97996 165034 98008
rect 213914 97996 213920 98008
rect 213972 97996 213978 98048
rect 258718 97996 258724 98048
rect 258776 98036 258782 98048
rect 307662 98036 307668 98048
rect 258776 98008 307668 98036
rect 258776 97996 258782 98008
rect 307662 97996 307668 98008
rect 307720 97996 307726 98048
rect 252462 97928 252468 97980
rect 252520 97968 252526 97980
rect 263042 97968 263048 97980
rect 252520 97940 263048 97968
rect 252520 97928 252526 97940
rect 263042 97928 263048 97940
rect 263100 97928 263106 97980
rect 2774 97724 2780 97776
rect 2832 97764 2838 97776
rect 4798 97764 4804 97776
rect 2832 97736 4804 97764
rect 2832 97724 2838 97736
rect 4798 97724 4804 97736
rect 4856 97724 4862 97776
rect 289354 96704 289360 96756
rect 289412 96744 289418 96756
rect 306926 96744 306932 96756
rect 289412 96716 306932 96744
rect 289412 96704 289418 96716
rect 306926 96704 306932 96716
rect 306984 96704 306990 96756
rect 210510 96636 210516 96688
rect 210568 96676 210574 96688
rect 213914 96676 213920 96688
rect 210568 96648 213920 96676
rect 210568 96636 210574 96648
rect 213914 96636 213920 96648
rect 213972 96636 213978 96688
rect 255958 96636 255964 96688
rect 256016 96676 256022 96688
rect 307662 96676 307668 96688
rect 256016 96648 307668 96676
rect 256016 96636 256022 96648
rect 307662 96636 307668 96648
rect 307720 96636 307726 96688
rect 308490 96568 308496 96620
rect 308548 96608 308554 96620
rect 321462 96608 321468 96620
rect 308548 96580 321468 96608
rect 308548 96568 308554 96580
rect 321462 96568 321468 96580
rect 321520 96568 321526 96620
rect 198182 95208 198188 95260
rect 198240 95248 198246 95260
rect 213914 95248 213920 95260
rect 198240 95220 213920 95248
rect 198240 95208 198246 95220
rect 213914 95208 213920 95220
rect 213972 95208 213978 95260
rect 249058 95208 249064 95260
rect 249116 95248 249122 95260
rect 307662 95248 307668 95260
rect 249116 95220 307668 95248
rect 249116 95208 249122 95220
rect 307662 95208 307668 95220
rect 307720 95208 307726 95260
rect 196618 95140 196624 95192
rect 196676 95180 196682 95192
rect 324314 95180 324320 95192
rect 196676 95152 324320 95180
rect 196676 95140 196682 95152
rect 324314 95140 324320 95152
rect 324372 95140 324378 95192
rect 308398 95072 308404 95124
rect 308456 95112 308462 95124
rect 324406 95112 324412 95124
rect 308456 95084 324412 95112
rect 308456 95072 308462 95084
rect 324406 95072 324412 95084
rect 324464 95072 324470 95124
rect 309778 95004 309784 95056
rect 309836 95044 309842 95056
rect 321370 95044 321376 95056
rect 309836 95016 321376 95044
rect 309836 95004 309842 95016
rect 321370 95004 321376 95016
rect 321428 95004 321434 95056
rect 122834 94460 122840 94512
rect 122892 94500 122898 94512
rect 214834 94500 214840 94512
rect 122892 94472 214840 94500
rect 122892 94460 122898 94472
rect 214834 94460 214840 94472
rect 214892 94460 214898 94512
rect 151630 94052 151636 94104
rect 151688 94092 151694 94104
rect 178678 94092 178684 94104
rect 151688 94064 178684 94092
rect 151688 94052 151694 94064
rect 178678 94052 178684 94064
rect 178736 94052 178742 94104
rect 129366 93984 129372 94036
rect 129424 94024 129430 94036
rect 166258 94024 166264 94036
rect 129424 93996 166264 94024
rect 129424 93984 129430 93996
rect 166258 93984 166264 93996
rect 166316 93984 166322 94036
rect 111978 93916 111984 93968
rect 112036 93956 112042 93968
rect 170490 93956 170496 93968
rect 112036 93928 170496 93956
rect 112036 93916 112042 93928
rect 170490 93916 170496 93928
rect 170548 93916 170554 93968
rect 113726 93848 113732 93900
rect 113784 93888 113790 93900
rect 172054 93888 172060 93900
rect 113784 93860 172060 93888
rect 113784 93848 113790 93860
rect 172054 93848 172060 93860
rect 172112 93848 172118 93900
rect 62022 93780 62028 93832
rect 62080 93820 62086 93832
rect 210602 93820 210608 93832
rect 62080 93792 210608 93820
rect 62080 93780 62086 93792
rect 210602 93780 210608 93792
rect 210660 93780 210666 93832
rect 216030 93780 216036 93832
rect 216088 93820 216094 93832
rect 321646 93820 321652 93832
rect 216088 93792 321652 93820
rect 216088 93780 216094 93792
rect 321646 93780 321652 93792
rect 321704 93780 321710 93832
rect 188338 93712 188344 93764
rect 188396 93752 188402 93764
rect 324498 93752 324504 93764
rect 188396 93724 324504 93752
rect 188396 93712 188402 93724
rect 324498 93712 324504 93724
rect 324556 93712 324562 93764
rect 191098 93644 191104 93696
rect 191156 93684 191162 93696
rect 321554 93684 321560 93696
rect 191156 93656 321560 93684
rect 191156 93644 191162 93656
rect 321554 93644 321560 93656
rect 321612 93644 321618 93696
rect 133138 93372 133144 93424
rect 133196 93412 133202 93424
rect 174538 93412 174544 93424
rect 133196 93384 174544 93412
rect 133196 93372 133202 93384
rect 174538 93372 174544 93384
rect 174596 93372 174602 93424
rect 118050 93304 118056 93356
rect 118108 93344 118114 93356
rect 170398 93344 170404 93356
rect 118108 93316 170404 93344
rect 118108 93304 118114 93316
rect 170398 93304 170404 93316
rect 170456 93304 170462 93356
rect 120626 93236 120632 93288
rect 120684 93276 120690 93288
rect 195330 93276 195336 93288
rect 120684 93248 195336 93276
rect 120684 93236 120690 93248
rect 195330 93236 195336 93248
rect 195388 93236 195394 93288
rect 107746 93168 107752 93220
rect 107804 93208 107810 93220
rect 186958 93208 186964 93220
rect 107804 93180 186964 93208
rect 107804 93168 107810 93180
rect 186958 93168 186964 93180
rect 187016 93168 187022 93220
rect 85666 93100 85672 93152
rect 85724 93140 85730 93152
rect 164970 93140 164976 93152
rect 85724 93112 164976 93140
rect 85724 93100 85730 93112
rect 164970 93100 164976 93112
rect 165028 93100 165034 93152
rect 115474 92420 115480 92472
rect 115532 92460 115538 92472
rect 204898 92460 204904 92472
rect 115532 92432 204904 92460
rect 115532 92420 115538 92432
rect 204898 92420 204904 92432
rect 204956 92420 204962 92472
rect 95050 92352 95056 92404
rect 95108 92392 95114 92404
rect 122834 92392 122840 92404
rect 95108 92364 122840 92392
rect 95108 92352 95114 92364
rect 122834 92352 122840 92364
rect 122892 92352 122898 92404
rect 125962 92352 125968 92404
rect 126020 92392 126026 92404
rect 206370 92392 206376 92404
rect 126020 92364 206376 92392
rect 126020 92352 126026 92364
rect 206370 92352 206376 92364
rect 206428 92352 206434 92404
rect 116762 92284 116768 92336
rect 116820 92324 116826 92336
rect 174722 92324 174728 92336
rect 116820 92296 174728 92324
rect 116820 92284 116826 92296
rect 174722 92284 174728 92296
rect 174780 92284 174786 92336
rect 151722 92216 151728 92268
rect 151780 92256 151786 92268
rect 197998 92256 198004 92268
rect 151780 92228 198004 92256
rect 151780 92216 151786 92228
rect 197998 92216 198004 92228
rect 198056 92216 198062 92268
rect 130746 92148 130752 92200
rect 130804 92188 130810 92200
rect 169018 92188 169024 92200
rect 130804 92160 169024 92188
rect 130804 92148 130810 92160
rect 169018 92148 169024 92160
rect 169076 92148 169082 92200
rect 152090 92080 152096 92132
rect 152148 92120 152154 92132
rect 173250 92120 173256 92132
rect 152148 92092 173256 92120
rect 152148 92080 152154 92092
rect 173250 92080 173256 92092
rect 173308 92080 173314 92132
rect 238018 91808 238024 91860
rect 238076 91848 238082 91860
rect 251174 91848 251180 91860
rect 238076 91820 251180 91848
rect 238076 91808 238082 91820
rect 251174 91808 251180 91820
rect 251232 91808 251238 91860
rect 206278 91740 206284 91792
rect 206336 91780 206342 91792
rect 307294 91780 307300 91792
rect 206336 91752 307300 91780
rect 206336 91740 206342 91752
rect 307294 91740 307300 91752
rect 307352 91740 307358 91792
rect 91646 91128 91652 91180
rect 91704 91168 91710 91180
rect 108298 91168 108304 91180
rect 91704 91140 108304 91168
rect 91704 91128 91710 91140
rect 108298 91128 108304 91140
rect 108356 91128 108362 91180
rect 85114 91060 85120 91112
rect 85172 91100 85178 91112
rect 128998 91100 129004 91112
rect 85172 91072 129004 91100
rect 85172 91060 85178 91072
rect 128998 91060 129004 91072
rect 129056 91060 129062 91112
rect 66070 90992 66076 91044
rect 66128 91032 66134 91044
rect 171962 91032 171968 91044
rect 66128 91004 171968 91032
rect 66128 90992 66134 91004
rect 171962 90992 171968 91004
rect 172020 90992 172026 91044
rect 120534 90924 120540 90976
rect 120592 90964 120598 90976
rect 209038 90964 209044 90976
rect 120592 90936 209044 90964
rect 120592 90924 120598 90936
rect 209038 90924 209044 90936
rect 209096 90924 209102 90976
rect 105998 90856 106004 90908
rect 106056 90896 106062 90908
rect 189718 90896 189724 90908
rect 106056 90868 189724 90896
rect 106056 90856 106062 90868
rect 189718 90856 189724 90868
rect 189776 90856 189782 90908
rect 110322 90788 110328 90840
rect 110380 90828 110386 90840
rect 176102 90828 176108 90840
rect 110380 90800 176108 90828
rect 110380 90788 110386 90800
rect 176102 90788 176108 90800
rect 176160 90788 176166 90840
rect 125502 90720 125508 90772
rect 125560 90760 125566 90772
rect 169110 90760 169116 90772
rect 125560 90732 169116 90760
rect 125560 90720 125566 90732
rect 169110 90720 169116 90732
rect 169168 90720 169174 90772
rect 136450 90652 136456 90704
rect 136508 90692 136514 90704
rect 167730 90692 167736 90704
rect 136508 90664 167736 90692
rect 136508 90652 136514 90664
rect 167730 90652 167736 90664
rect 167788 90652 167794 90704
rect 177298 90312 177304 90364
rect 177356 90352 177362 90364
rect 307202 90352 307208 90364
rect 177356 90324 307208 90352
rect 177356 90312 177362 90324
rect 307202 90312 307208 90324
rect 307260 90312 307266 90364
rect 64782 89632 64788 89684
rect 64840 89672 64846 89684
rect 216214 89672 216220 89684
rect 64840 89644 216220 89672
rect 64840 89632 64846 89644
rect 216214 89632 216220 89644
rect 216272 89632 216278 89684
rect 90634 89564 90640 89616
rect 90692 89604 90698 89616
rect 199470 89604 199476 89616
rect 90692 89576 199476 89604
rect 90692 89564 90698 89576
rect 199470 89564 199476 89576
rect 199528 89564 199534 89616
rect 102686 89496 102692 89548
rect 102744 89536 102750 89548
rect 211890 89536 211896 89548
rect 102744 89508 211896 89536
rect 102744 89496 102750 89508
rect 211890 89496 211896 89508
rect 211948 89496 211954 89548
rect 100018 89428 100024 89480
rect 100076 89468 100082 89480
rect 192478 89468 192484 89480
rect 100076 89440 192484 89468
rect 100076 89428 100082 89440
rect 192478 89428 192484 89440
rect 192536 89428 192542 89480
rect 115382 89360 115388 89412
rect 115440 89400 115446 89412
rect 178862 89400 178868 89412
rect 115440 89372 178868 89400
rect 115440 89360 115446 89372
rect 178862 89360 178868 89372
rect 178920 89360 178926 89412
rect 151262 89292 151268 89344
rect 151320 89332 151326 89344
rect 213178 89332 213184 89344
rect 151320 89304 213184 89332
rect 151320 89292 151326 89304
rect 213178 89292 213184 89304
rect 213236 89292 213242 89344
rect 215938 88952 215944 89004
rect 215996 88992 216002 89004
rect 307110 88992 307116 89004
rect 215996 88964 307116 88992
rect 215996 88952 216002 88964
rect 307110 88952 307116 88964
rect 307168 88952 307174 89004
rect 67634 88272 67640 88324
rect 67692 88312 67698 88324
rect 214926 88312 214932 88324
rect 67692 88284 214932 88312
rect 67692 88272 67698 88284
rect 214926 88272 214932 88284
rect 214984 88272 214990 88324
rect 67450 88204 67456 88256
rect 67508 88244 67514 88256
rect 214558 88244 214564 88256
rect 67508 88216 214564 88244
rect 67508 88204 67514 88216
rect 214558 88204 214564 88216
rect 214616 88204 214622 88256
rect 126514 88136 126520 88188
rect 126572 88176 126578 88188
rect 191190 88176 191196 88188
rect 126572 88148 191196 88176
rect 126572 88136 126578 88148
rect 191190 88136 191196 88148
rect 191248 88136 191254 88188
rect 111242 88068 111248 88120
rect 111300 88108 111306 88120
rect 167822 88108 167828 88120
rect 111300 88080 167828 88108
rect 111300 88068 111306 88080
rect 167822 88068 167828 88080
rect 167880 88068 167886 88120
rect 117130 88000 117136 88052
rect 117188 88040 117194 88052
rect 170674 88040 170680 88052
rect 117188 88012 170680 88040
rect 117188 88000 117194 88012
rect 170674 88000 170680 88012
rect 170732 88000 170738 88052
rect 123478 87932 123484 87984
rect 123536 87972 123542 87984
rect 177390 87972 177396 87984
rect 123536 87944 177396 87972
rect 123536 87932 123542 87944
rect 177390 87932 177396 87944
rect 177448 87932 177454 87984
rect 101858 86912 101864 86964
rect 101916 86952 101922 86964
rect 204990 86952 204996 86964
rect 101916 86924 204996 86952
rect 101916 86912 101922 86924
rect 204990 86912 204996 86924
rect 205048 86912 205054 86964
rect 88058 86844 88064 86896
rect 88116 86884 88122 86896
rect 166534 86884 166540 86896
rect 88116 86856 166540 86884
rect 88116 86844 88122 86856
rect 166534 86844 166540 86856
rect 166592 86844 166598 86896
rect 134610 86776 134616 86828
rect 134668 86816 134674 86828
rect 210418 86816 210424 86828
rect 134668 86788 210424 86816
rect 134668 86776 134674 86788
rect 210418 86776 210424 86788
rect 210476 86776 210482 86828
rect 109586 86708 109592 86760
rect 109644 86748 109650 86760
rect 177482 86748 177488 86760
rect 109644 86720 177488 86748
rect 109644 86708 109650 86720
rect 177482 86708 177488 86720
rect 177540 86708 177546 86760
rect 112346 86640 112352 86692
rect 112404 86680 112410 86692
rect 167914 86680 167920 86692
rect 112404 86652 167920 86680
rect 112404 86640 112410 86652
rect 167914 86640 167920 86652
rect 167972 86640 167978 86692
rect 124122 86572 124128 86624
rect 124180 86612 124186 86624
rect 170582 86612 170588 86624
rect 124180 86584 170588 86612
rect 124180 86572 124186 86584
rect 170582 86572 170588 86584
rect 170640 86572 170646 86624
rect 3510 85484 3516 85536
rect 3568 85524 3574 85536
rect 22738 85524 22744 85536
rect 3568 85496 22744 85524
rect 3568 85484 3574 85496
rect 22738 85484 22744 85496
rect 22796 85484 22802 85536
rect 67358 85484 67364 85536
rect 67416 85524 67422 85536
rect 210510 85524 210516 85536
rect 67416 85496 210516 85524
rect 67416 85484 67422 85496
rect 210510 85484 210516 85496
rect 210568 85484 210574 85536
rect 111426 85416 111432 85468
rect 111484 85456 111490 85468
rect 213362 85456 213368 85468
rect 111484 85428 213368 85456
rect 111484 85416 111490 85428
rect 213362 85416 213368 85428
rect 213420 85416 213426 85468
rect 104250 85348 104256 85400
rect 104308 85388 104314 85400
rect 198090 85388 198096 85400
rect 104308 85360 198096 85388
rect 104308 85348 104314 85360
rect 198090 85348 198096 85360
rect 198148 85348 198154 85400
rect 100570 85280 100576 85332
rect 100628 85320 100634 85332
rect 169202 85320 169208 85332
rect 100628 85292 169208 85320
rect 100628 85280 100634 85292
rect 169202 85280 169208 85292
rect 169260 85280 169266 85332
rect 122834 85212 122840 85264
rect 122892 85252 122898 85264
rect 180058 85252 180064 85264
rect 122892 85224 180064 85252
rect 122892 85212 122898 85224
rect 180058 85212 180064 85224
rect 180116 85212 180122 85264
rect 132402 85144 132408 85196
rect 132460 85184 132466 85196
rect 173158 85184 173164 85196
rect 132460 85156 173164 85184
rect 132460 85144 132466 85156
rect 173158 85144 173164 85156
rect 173216 85144 173222 85196
rect 104802 84124 104808 84176
rect 104860 84164 104866 84176
rect 207658 84164 207664 84176
rect 104860 84136 207664 84164
rect 104860 84124 104866 84136
rect 207658 84124 207664 84136
rect 207716 84124 207722 84176
rect 118602 84056 118608 84108
rect 118660 84096 118666 84108
rect 202230 84096 202236 84108
rect 118660 84068 202236 84096
rect 118660 84056 118666 84068
rect 202230 84056 202236 84068
rect 202288 84056 202294 84108
rect 86862 83988 86868 84040
rect 86920 84028 86926 84040
rect 166442 84028 166448 84040
rect 86920 84000 166448 84028
rect 86920 83988 86926 84000
rect 166442 83988 166448 84000
rect 166500 83988 166506 84040
rect 96522 83920 96528 83972
rect 96580 83960 96586 83972
rect 174630 83960 174636 83972
rect 96580 83932 174636 83960
rect 96580 83920 96586 83932
rect 174630 83920 174636 83932
rect 174688 83920 174694 83972
rect 106182 83852 106188 83904
rect 106240 83892 106246 83904
rect 180150 83892 180156 83904
rect 106240 83864 180156 83892
rect 106240 83852 106246 83864
rect 180150 83852 180156 83864
rect 180208 83852 180214 83904
rect 122650 83784 122656 83836
rect 122708 83824 122714 83836
rect 171778 83824 171784 83836
rect 122708 83796 171784 83824
rect 122708 83784 122714 83796
rect 171778 83784 171784 83796
rect 171836 83784 171842 83836
rect 122742 82764 122748 82816
rect 122800 82804 122806 82816
rect 211798 82804 211804 82816
rect 122800 82776 211804 82804
rect 122800 82764 122806 82776
rect 211798 82764 211804 82776
rect 211856 82764 211862 82816
rect 89622 82696 89628 82748
rect 89680 82736 89686 82748
rect 166350 82736 166356 82748
rect 89680 82708 166356 82736
rect 89680 82696 89686 82708
rect 166350 82696 166356 82708
rect 166408 82696 166414 82748
rect 99098 82628 99104 82680
rect 99156 82668 99162 82680
rect 173434 82668 173440 82680
rect 99156 82640 173440 82668
rect 99156 82628 99162 82640
rect 173434 82628 173440 82640
rect 173492 82628 173498 82680
rect 110138 82560 110144 82612
rect 110196 82600 110202 82612
rect 181438 82600 181444 82612
rect 110196 82572 181444 82600
rect 110196 82560 110202 82572
rect 181438 82560 181444 82572
rect 181496 82560 181502 82612
rect 101950 82492 101956 82544
rect 102008 82532 102014 82544
rect 171870 82532 171876 82544
rect 102008 82504 171876 82532
rect 102008 82492 102014 82504
rect 171870 82492 171876 82504
rect 171928 82492 171934 82544
rect 125410 82424 125416 82476
rect 125468 82464 125474 82476
rect 167638 82464 167644 82476
rect 125468 82436 167644 82464
rect 125468 82424 125474 82436
rect 167638 82424 167644 82436
rect 167696 82424 167702 82476
rect 108298 81336 108304 81388
rect 108356 81376 108362 81388
rect 214650 81376 214656 81388
rect 108356 81348 214656 81376
rect 108356 81336 108362 81348
rect 214650 81336 214656 81348
rect 214708 81336 214714 81388
rect 93762 81268 93768 81320
rect 93820 81308 93826 81320
rect 169294 81308 169300 81320
rect 93820 81280 169300 81308
rect 93820 81268 93826 81280
rect 169294 81268 169300 81280
rect 169352 81268 169358 81320
rect 128262 81200 128268 81252
rect 128320 81240 128326 81252
rect 202138 81240 202144 81252
rect 128320 81212 202144 81240
rect 128320 81200 128326 81212
rect 202138 81200 202144 81212
rect 202196 81200 202202 81252
rect 107470 81132 107476 81184
rect 107528 81172 107534 81184
rect 173342 81172 173348 81184
rect 107528 81144 173348 81172
rect 107528 81132 107534 81144
rect 173342 81132 173348 81144
rect 173400 81132 173406 81184
rect 115842 79976 115848 80028
rect 115900 80016 115906 80028
rect 213270 80016 213276 80028
rect 115900 79988 213276 80016
rect 115900 79976 115906 79988
rect 213270 79976 213276 79988
rect 213328 79976 213334 80028
rect 108942 79908 108948 79960
rect 109000 79948 109006 79960
rect 196710 79948 196716 79960
rect 109000 79920 196716 79948
rect 109000 79908 109006 79920
rect 196710 79908 196716 79920
rect 196768 79908 196774 79960
rect 95142 79840 95148 79892
rect 95200 79880 95206 79892
rect 177666 79880 177672 79892
rect 95200 79852 177672 79880
rect 95200 79840 95206 79852
rect 177666 79840 177672 79852
rect 177724 79840 177730 79892
rect 114462 79772 114468 79824
rect 114520 79812 114526 79824
rect 195238 79812 195244 79824
rect 114520 79784 195244 79812
rect 114520 79772 114526 79784
rect 195238 79772 195244 79784
rect 195296 79772 195302 79824
rect 97902 78616 97908 78668
rect 97960 78656 97966 78668
rect 209130 78656 209136 78668
rect 97960 78628 209136 78656
rect 97960 78616 97966 78628
rect 209130 78616 209136 78628
rect 209188 78616 209194 78668
rect 128998 78548 129004 78600
rect 129056 78588 129062 78600
rect 216122 78588 216128 78600
rect 129056 78560 216128 78588
rect 129056 78548 129062 78560
rect 216122 78548 216128 78560
rect 216180 78548 216186 78600
rect 102042 78480 102048 78532
rect 102100 78520 102106 78532
rect 178770 78520 178776 78532
rect 102100 78492 178776 78520
rect 102100 78480 102106 78492
rect 178770 78480 178776 78492
rect 178828 78480 178834 78532
rect 119982 78412 119988 78464
rect 120040 78452 120046 78464
rect 182818 78452 182824 78464
rect 120040 78424 182824 78452
rect 120040 78412 120046 78424
rect 182818 78412 182824 78424
rect 182876 78412 182882 78464
rect 75822 77188 75828 77240
rect 75880 77228 75886 77240
rect 198182 77228 198188 77240
rect 75880 77200 198188 77228
rect 75880 77188 75886 77200
rect 198182 77188 198188 77200
rect 198240 77188 198246 77240
rect 124214 76576 124220 76628
rect 124272 76616 124278 76628
rect 279510 76616 279516 76628
rect 124272 76588 279516 76616
rect 124272 76576 124278 76588
rect 279510 76576 279516 76588
rect 279568 76576 279574 76628
rect 82814 76508 82820 76560
rect 82872 76548 82878 76560
rect 292206 76548 292212 76560
rect 82872 76520 292212 76548
rect 82872 76508 82878 76520
rect 292206 76508 292212 76520
rect 292264 76508 292270 76560
rect 107562 75828 107568 75880
rect 107620 75868 107626 75880
rect 176010 75868 176016 75880
rect 107620 75840 176016 75868
rect 107620 75828 107626 75840
rect 176010 75828 176016 75840
rect 176068 75828 176074 75880
rect 115934 75216 115940 75268
rect 115992 75256 115998 75268
rect 303062 75256 303068 75268
rect 115992 75228 303068 75256
rect 115992 75216 115998 75228
rect 303062 75216 303068 75228
rect 303120 75216 303126 75268
rect 23474 75148 23480 75200
rect 23532 75188 23538 75200
rect 272518 75188 272524 75200
rect 23532 75160 272524 75188
rect 23532 75148 23538 75160
rect 272518 75148 272524 75160
rect 272576 75148 272582 75200
rect 93854 73856 93860 73908
rect 93912 73896 93918 73908
rect 306006 73896 306012 73908
rect 93912 73868 306012 73896
rect 93912 73856 93918 73868
rect 306006 73856 306012 73868
rect 306064 73856 306070 73908
rect 56594 73788 56600 73840
rect 56652 73828 56658 73840
rect 294782 73828 294788 73840
rect 56652 73800 294788 73828
rect 56652 73788 56658 73800
rect 294782 73788 294788 73800
rect 294840 73788 294846 73840
rect 118694 72496 118700 72548
rect 118752 72536 118758 72548
rect 298922 72536 298928 72548
rect 118752 72508 298928 72536
rect 118752 72496 118758 72508
rect 298922 72496 298928 72508
rect 298980 72496 298986 72548
rect 64874 72428 64880 72480
rect 64932 72468 64938 72480
rect 300486 72468 300492 72480
rect 64932 72440 300492 72468
rect 64932 72428 64938 72440
rect 300486 72428 300492 72440
rect 300544 72428 300550 72480
rect 3510 71680 3516 71732
rect 3568 71720 3574 71732
rect 53098 71720 53104 71732
rect 3568 71692 53104 71720
rect 3568 71680 3574 71692
rect 53098 71680 53104 71692
rect 53156 71680 53162 71732
rect 103514 71068 103520 71120
rect 103572 71108 103578 71120
rect 304534 71108 304540 71120
rect 103572 71080 304540 71108
rect 103572 71068 103578 71080
rect 304534 71068 304540 71080
rect 304592 71068 304598 71120
rect 52454 71000 52460 71052
rect 52512 71040 52518 71052
rect 296254 71040 296260 71052
rect 52512 71012 296260 71040
rect 52512 71000 52518 71012
rect 296254 71000 296260 71012
rect 296312 71000 296318 71052
rect 9674 69640 9680 69692
rect 9732 69680 9738 69692
rect 286502 69680 286508 69692
rect 9732 69652 286508 69680
rect 9732 69640 9738 69652
rect 286502 69640 286508 69652
rect 286560 69640 286566 69692
rect 110414 68348 110420 68400
rect 110472 68388 110478 68400
rect 303154 68388 303160 68400
rect 110472 68360 303160 68388
rect 110472 68348 110478 68360
rect 303154 68348 303160 68360
rect 303212 68348 303218 68400
rect 44174 68280 44180 68332
rect 44232 68320 44238 68332
rect 267182 68320 267188 68332
rect 44232 68292 267188 68320
rect 44232 68280 44238 68292
rect 267182 68280 267188 68292
rect 267240 68280 267246 68332
rect 114554 66920 114560 66972
rect 114612 66960 114618 66972
rect 300210 66960 300216 66972
rect 114612 66932 300216 66960
rect 114612 66920 114618 66932
rect 300210 66920 300216 66932
rect 300268 66920 300274 66972
rect 34514 66852 34520 66904
rect 34572 66892 34578 66904
rect 293402 66892 293408 66904
rect 34572 66864 293408 66892
rect 34572 66852 34578 66864
rect 293402 66852 293408 66864
rect 293460 66852 293466 66904
rect 121454 65560 121460 65612
rect 121512 65600 121518 65612
rect 253198 65600 253204 65612
rect 121512 65572 253204 65600
rect 121512 65560 121518 65572
rect 253198 65560 253204 65572
rect 253256 65560 253262 65612
rect 30374 65492 30380 65544
rect 30432 65532 30438 65544
rect 287882 65532 287888 65544
rect 30432 65504 287888 65532
rect 30432 65492 30438 65504
rect 287882 65492 287888 65504
rect 287940 65492 287946 65544
rect 69014 64200 69020 64252
rect 69072 64240 69078 64252
rect 305822 64240 305828 64252
rect 69072 64212 305828 64240
rect 69072 64200 69078 64212
rect 305822 64200 305828 64212
rect 305880 64200 305886 64252
rect 28994 64132 29000 64184
rect 29052 64172 29058 64184
rect 300394 64172 300400 64184
rect 29052 64144 300400 64172
rect 29052 64132 29058 64144
rect 300394 64132 300400 64144
rect 300452 64132 300458 64184
rect 71774 62772 71780 62824
rect 71832 62812 71838 62824
rect 268470 62812 268476 62824
rect 71832 62784 268476 62812
rect 71832 62772 71838 62784
rect 268470 62772 268476 62784
rect 268528 62772 268534 62824
rect 97994 61344 98000 61396
rect 98052 61384 98058 61396
rect 282362 61384 282368 61396
rect 98052 61356 282368 61384
rect 98052 61344 98058 61356
rect 282362 61344 282368 61356
rect 282420 61344 282426 61396
rect 184198 60664 184204 60716
rect 184256 60704 184262 60716
rect 580166 60704 580172 60716
rect 184256 60676 580172 60704
rect 184256 60664 184262 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 4154 59984 4160 60036
rect 4212 60024 4218 60036
rect 249058 60024 249064 60036
rect 4212 59996 249064 60024
rect 4212 59984 4218 59996
rect 249058 59984 249064 59996
rect 249116 59984 249122 60036
rect 70394 58692 70400 58744
rect 70452 58732 70458 58744
rect 290550 58732 290556 58744
rect 70452 58704 290556 58732
rect 70452 58692 70458 58704
rect 290550 58692 290556 58704
rect 290608 58692 290614 58744
rect 33134 58624 33140 58676
rect 33192 58664 33198 58676
rect 299014 58664 299020 58676
rect 33192 58636 299020 58664
rect 33192 58624 33198 58636
rect 299014 58624 299020 58636
rect 299072 58624 299078 58676
rect 85574 57196 85580 57248
rect 85632 57236 85638 57248
rect 291930 57236 291936 57248
rect 85632 57208 291936 57236
rect 85632 57196 85638 57208
rect 291930 57196 291936 57208
rect 291988 57196 291994 57248
rect 45554 55904 45560 55956
rect 45612 55944 45618 55956
rect 273990 55944 273996 55956
rect 45612 55916 273996 55944
rect 45612 55904 45618 55916
rect 273990 55904 273996 55916
rect 274048 55904 274054 55956
rect 73154 55836 73160 55888
rect 73212 55876 73218 55888
rect 301682 55876 301688 55888
rect 73212 55848 301688 55876
rect 73212 55836 73218 55848
rect 301682 55836 301688 55848
rect 301740 55836 301746 55888
rect 86954 53116 86960 53168
rect 87012 53156 87018 53168
rect 289262 53156 289268 53168
rect 87012 53128 289268 53156
rect 87012 53116 87018 53128
rect 289262 53116 289268 53128
rect 289320 53116 289326 53168
rect 27614 53048 27620 53100
rect 27672 53088 27678 53100
rect 271230 53088 271236 53100
rect 27672 53060 271236 53088
rect 27672 53048 27678 53060
rect 271230 53048 271236 53060
rect 271288 53048 271294 53100
rect 91094 51756 91100 51808
rect 91152 51796 91158 51808
rect 297542 51796 297548 51808
rect 91152 51768 297548 51796
rect 91152 51756 91158 51768
rect 297542 51756 297548 51768
rect 297600 51756 297606 51808
rect 19334 51688 19340 51740
rect 19392 51728 19398 51740
rect 289170 51728 289176 51740
rect 19392 51700 289176 51728
rect 19392 51688 19398 51700
rect 289170 51688 289176 51700
rect 289228 51688 289234 51740
rect 104894 50396 104900 50448
rect 104952 50436 104958 50448
rect 292022 50436 292028 50448
rect 104952 50408 292028 50436
rect 104952 50396 104958 50408
rect 292022 50396 292028 50408
rect 292080 50396 292086 50448
rect 81434 50328 81440 50380
rect 81492 50368 81498 50380
rect 276750 50368 276756 50380
rect 81492 50340 276756 50368
rect 81492 50328 81498 50340
rect 276750 50328 276756 50340
rect 276808 50328 276814 50380
rect 102134 49036 102140 49088
rect 102192 49076 102198 49088
rect 304350 49076 304356 49088
rect 102192 49048 304356 49076
rect 102192 49036 102198 49048
rect 304350 49036 304356 49048
rect 304408 49036 304414 49088
rect 60734 48968 60740 49020
rect 60792 49008 60798 49020
rect 271138 49008 271144 49020
rect 60792 48980 271144 49008
rect 60792 48968 60798 48980
rect 271138 48968 271144 48980
rect 271196 48968 271202 49020
rect 88334 47540 88340 47592
rect 88392 47580 88398 47592
rect 278130 47580 278136 47592
rect 88392 47552 278136 47580
rect 88392 47540 88398 47552
rect 278130 47540 278136 47552
rect 278188 47540 278194 47592
rect 14 46860 20 46912
rect 72 46900 78 46912
rect 1302 46900 1308 46912
rect 72 46872 1308 46900
rect 72 46860 78 46872
rect 1302 46860 1308 46872
rect 1360 46900 1366 46912
rect 249150 46900 249156 46912
rect 1360 46872 249156 46900
rect 1360 46860 1366 46872
rect 249150 46860 249156 46872
rect 249208 46860 249214 46912
rect 122834 46180 122840 46232
rect 122892 46220 122898 46232
rect 300118 46220 300124 46232
rect 122892 46192 300124 46220
rect 122892 46180 122898 46192
rect 300118 46180 300124 46192
rect 300176 46180 300182 46232
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 15838 45540 15844 45552
rect 3476 45512 15844 45540
rect 3476 45500 3482 45512
rect 15838 45500 15844 45512
rect 15896 45500 15902 45552
rect 93946 44888 93952 44940
rect 94004 44928 94010 44940
rect 286410 44928 286416 44940
rect 94004 44900 286416 44928
rect 94004 44888 94010 44900
rect 286410 44888 286416 44900
rect 286468 44888 286474 44940
rect 13814 44820 13820 44872
rect 13872 44860 13878 44872
rect 273898 44860 273904 44872
rect 13872 44832 273904 44860
rect 13872 44820 13878 44832
rect 273898 44820 273904 44832
rect 273956 44820 273962 44872
rect 84194 43460 84200 43512
rect 84252 43500 84258 43512
rect 269758 43500 269764 43512
rect 84252 43472 269764 43500
rect 84252 43460 84258 43472
rect 269758 43460 269764 43472
rect 269816 43460 269822 43512
rect 95234 43392 95240 43444
rect 95292 43432 95298 43444
rect 287698 43432 287704 43444
rect 95292 43404 287704 43432
rect 95292 43392 95298 43404
rect 287698 43392 287704 43404
rect 287756 43392 287762 43444
rect 80054 42100 80060 42152
rect 80112 42140 80118 42152
rect 290458 42140 290464 42152
rect 80112 42112 290464 42140
rect 80112 42100 80118 42112
rect 290458 42100 290464 42112
rect 290516 42100 290522 42152
rect 35986 42032 35992 42084
rect 36044 42072 36050 42084
rect 301590 42072 301596 42084
rect 36044 42044 301596 42072
rect 36044 42032 36050 42044
rect 301590 42032 301596 42044
rect 301648 42032 301654 42084
rect 77294 40740 77300 40792
rect 77352 40780 77358 40792
rect 291838 40780 291844 40792
rect 77352 40752 291844 40780
rect 77352 40740 77358 40752
rect 291838 40740 291844 40752
rect 291896 40740 291902 40792
rect 42794 40672 42800 40724
rect 42852 40712 42858 40724
rect 285122 40712 285128 40724
rect 42852 40684 285128 40712
rect 42852 40672 42858 40684
rect 285122 40672 285128 40684
rect 285180 40672 285186 40724
rect 57974 39380 57980 39432
rect 58032 39420 58038 39432
rect 267090 39420 267096 39432
rect 58032 39392 267096 39420
rect 58032 39380 58038 39392
rect 267090 39380 267096 39392
rect 267148 39380 267154 39432
rect 66254 39312 66260 39364
rect 66312 39352 66318 39364
rect 298830 39352 298836 39364
rect 66312 39324 298836 39352
rect 66312 39312 66318 39324
rect 298830 39312 298836 39324
rect 298888 39312 298894 39364
rect 99374 37952 99380 38004
rect 99432 37992 99438 38004
rect 283558 37992 283564 38004
rect 99432 37964 283564 37992
rect 99432 37952 99438 37964
rect 283558 37952 283564 37964
rect 283616 37952 283622 38004
rect 24854 37884 24860 37936
rect 24912 37924 24918 37936
rect 307018 37924 307024 37936
rect 24912 37896 307024 37924
rect 24912 37884 24918 37896
rect 307018 37884 307024 37896
rect 307076 37884 307082 37936
rect 92474 36592 92480 36644
rect 92532 36632 92538 36644
rect 302878 36632 302884 36644
rect 92532 36604 302884 36632
rect 92532 36592 92538 36604
rect 302878 36592 302884 36604
rect 302936 36592 302942 36644
rect 16574 36524 16580 36576
rect 16632 36564 16638 36576
rect 290642 36564 290648 36576
rect 16632 36536 290648 36564
rect 16632 36524 16638 36536
rect 290642 36524 290648 36536
rect 290700 36524 290706 36576
rect 40034 35232 40040 35284
rect 40092 35272 40098 35284
rect 269850 35272 269856 35284
rect 40092 35244 269856 35272
rect 40092 35232 40098 35244
rect 269850 35232 269856 35244
rect 269908 35232 269914 35284
rect 52546 35164 52552 35216
rect 52604 35204 52610 35216
rect 293310 35204 293316 35216
rect 52604 35176 293316 35204
rect 52604 35164 52610 35176
rect 293310 35164 293316 35176
rect 293368 35164 293374 35216
rect 106274 33804 106280 33856
rect 106332 33844 106338 33856
rect 293218 33844 293224 33856
rect 106332 33816 293224 33844
rect 106332 33804 106338 33816
rect 293218 33804 293224 33816
rect 293276 33804 293282 33856
rect 48314 33736 48320 33788
rect 48372 33776 48378 33788
rect 296162 33776 296168 33788
rect 48372 33748 296168 33776
rect 48372 33736 48378 33748
rect 296162 33736 296168 33748
rect 296220 33736 296226 33788
rect 3142 33056 3148 33108
rect 3200 33096 3206 33108
rect 32398 33096 32404 33108
rect 3200 33068 32404 33096
rect 3200 33056 3206 33068
rect 32398 33056 32404 33068
rect 32456 33056 32462 33108
rect 2774 31016 2780 31068
rect 2832 31056 2838 31068
rect 289354 31056 289360 31068
rect 2832 31028 289360 31056
rect 2832 31016 2838 31028
rect 289354 31016 289360 31028
rect 289412 31016 289418 31068
rect 44266 29588 44272 29640
rect 44324 29628 44330 29640
rect 294690 29628 294696 29640
rect 44324 29600 294696 29628
rect 44324 29588 44330 29600
rect 294690 29588 294696 29600
rect 294748 29588 294754 29640
rect 75914 28296 75920 28348
rect 75972 28336 75978 28348
rect 305730 28336 305736 28348
rect 75972 28308 305736 28336
rect 75972 28296 75978 28308
rect 305730 28296 305736 28308
rect 305788 28296 305794 28348
rect 26234 28228 26240 28280
rect 26292 28268 26298 28280
rect 283650 28268 283656 28280
rect 26292 28240 283656 28268
rect 26292 28228 26298 28240
rect 283650 28228 283656 28240
rect 283708 28228 283714 28280
rect 96614 26936 96620 26988
rect 96672 26976 96678 26988
rect 262858 26976 262864 26988
rect 96672 26948 262864 26976
rect 96672 26936 96678 26948
rect 262858 26936 262864 26948
rect 262916 26936 262922 26988
rect 20714 26868 20720 26920
rect 20772 26908 20778 26920
rect 297450 26908 297456 26920
rect 20772 26880 297456 26908
rect 20772 26868 20778 26880
rect 297450 26868 297456 26880
rect 297508 26868 297514 26920
rect 118786 25576 118792 25628
rect 118844 25616 118850 25628
rect 301498 25616 301504 25628
rect 118844 25588 301504 25616
rect 118844 25576 118850 25588
rect 301498 25576 301504 25588
rect 301556 25576 301562 25628
rect 37274 25508 37280 25560
rect 37332 25548 37338 25560
rect 264238 25548 264244 25560
rect 37332 25520 264244 25548
rect 37332 25508 37338 25520
rect 264238 25508 264244 25520
rect 264296 25508 264302 25560
rect 107654 24148 107660 24200
rect 107712 24188 107718 24200
rect 305638 24188 305644 24200
rect 107712 24160 305644 24188
rect 107712 24148 107718 24160
rect 305638 24148 305644 24160
rect 305696 24148 305702 24200
rect 41414 24080 41420 24132
rect 41472 24120 41478 24132
rect 280890 24120 280896 24132
rect 41472 24092 280896 24120
rect 41472 24080 41478 24092
rect 280890 24080 280896 24092
rect 280948 24080 280954 24132
rect 100754 22788 100760 22840
rect 100812 22828 100818 22840
rect 287790 22828 287796 22840
rect 100812 22800 287796 22828
rect 100812 22788 100818 22800
rect 287790 22788 287796 22800
rect 287848 22788 287854 22840
rect 63494 22720 63500 22772
rect 63552 22760 63558 22772
rect 278038 22760 278044 22772
rect 63552 22732 278044 22760
rect 63552 22720 63558 22732
rect 278038 22720 278044 22732
rect 278096 22720 278102 22772
rect 85666 21428 85672 21480
rect 85724 21468 85730 21480
rect 302970 21468 302976 21480
rect 85724 21440 302976 21468
rect 85724 21428 85730 21440
rect 302970 21428 302976 21440
rect 303028 21428 303034 21480
rect 31754 21360 31760 21412
rect 31812 21400 31818 21412
rect 296070 21400 296076 21412
rect 31812 21372 296076 21400
rect 31812 21360 31818 21372
rect 296070 21360 296076 21372
rect 296128 21360 296134 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 11698 20652 11704 20664
rect 3476 20624 11704 20652
rect 3476 20612 3482 20624
rect 11698 20612 11704 20624
rect 11756 20612 11762 20664
rect 17954 19932 17960 19984
rect 18012 19972 18018 19984
rect 294598 19972 294604 19984
rect 18012 19944 294604 19972
rect 18012 19932 18018 19944
rect 294598 19932 294604 19944
rect 294656 19932 294662 19984
rect 89714 18572 89720 18624
rect 89772 18612 89778 18624
rect 282270 18612 282276 18624
rect 89772 18584 282276 18612
rect 89772 18572 89778 18584
rect 282270 18572 282276 18584
rect 282328 18572 282334 18624
rect 78674 17280 78680 17332
rect 78732 17320 78738 17332
rect 304258 17320 304264 17332
rect 78732 17292 304264 17320
rect 78732 17280 78738 17292
rect 304258 17280 304264 17292
rect 304316 17280 304322 17332
rect 38654 17212 38660 17264
rect 38712 17252 38718 17264
rect 276658 17252 276664 17264
rect 38712 17224 276664 17252
rect 38712 17212 38718 17224
rect 276658 17212 276664 17224
rect 276716 17212 276722 17264
rect 69106 15920 69112 15972
rect 69164 15960 69170 15972
rect 298738 15960 298744 15972
rect 69164 15932 298744 15960
rect 69164 15920 69170 15932
rect 298738 15920 298744 15932
rect 298796 15920 298802 15972
rect 11146 15852 11152 15904
rect 11204 15892 11210 15904
rect 255958 15892 255964 15904
rect 11204 15864 255964 15892
rect 11204 15852 11210 15864
rect 255958 15852 255964 15864
rect 256016 15852 256022 15904
rect 61562 14492 61568 14544
rect 61620 14532 61626 14544
rect 285030 14532 285036 14544
rect 61620 14504 285036 14532
rect 61620 14492 61626 14504
rect 285030 14492 285036 14504
rect 285088 14492 285094 14544
rect 20162 14424 20168 14476
rect 20220 14464 20226 14476
rect 258718 14464 258724 14476
rect 20220 14436 258724 14464
rect 20220 14424 20226 14436
rect 258718 14424 258724 14436
rect 258776 14424 258782 14476
rect 3418 13132 3424 13184
rect 3476 13172 3482 13184
rect 51718 13172 51724 13184
rect 3476 13144 51724 13172
rect 3476 13132 3482 13144
rect 51718 13132 51724 13144
rect 51776 13132 51782 13184
rect 51074 13064 51080 13116
rect 51132 13104 51138 13116
rect 279418 13104 279424 13116
rect 51132 13076 279424 13104
rect 51132 13064 51138 13076
rect 279418 13064 279424 13076
rect 279476 13064 279482 13116
rect 120626 11772 120632 11824
rect 120684 11812 120690 11824
rect 250438 11812 250444 11824
rect 120684 11784 250444 11812
rect 120684 11772 120690 11784
rect 250438 11772 250444 11784
rect 250496 11772 250502 11824
rect 7650 11704 7656 11756
rect 7708 11744 7714 11756
rect 286318 11744 286324 11756
rect 7708 11716 286324 11744
rect 7708 11704 7714 11716
rect 286318 11704 286324 11716
rect 286376 11704 286382 11756
rect 117314 10344 117320 10396
rect 117372 10384 117378 10396
rect 266998 10384 267004 10396
rect 117372 10356 267004 10384
rect 117372 10344 117378 10356
rect 266998 10344 267004 10356
rect 267056 10344 267062 10396
rect 2866 10276 2872 10328
rect 2924 10316 2930 10328
rect 289078 10316 289084 10328
rect 2924 10288 289084 10316
rect 2924 10276 2930 10288
rect 289078 10276 289084 10288
rect 289136 10276 289142 10328
rect 7466 9596 7472 9648
rect 7524 9636 7530 9648
rect 8202 9636 8208 9648
rect 7524 9608 8208 9636
rect 7524 9596 7530 9608
rect 8202 9596 8208 9608
rect 8260 9636 8266 9648
rect 251174 9636 251180 9648
rect 8260 9608 251180 9636
rect 8260 9596 8266 9608
rect 251174 9596 251180 9608
rect 251232 9596 251238 9648
rect 74994 8916 75000 8968
rect 75052 8956 75058 8968
rect 282178 8956 282184 8968
rect 75052 8928 282184 8956
rect 75052 8916 75058 8928
rect 282178 8916 282184 8928
rect 282236 8916 282242 8968
rect 1670 8304 1676 8356
rect 1728 8344 1734 8356
rect 7466 8344 7472 8356
rect 1728 8316 7472 8344
rect 1728 8304 1734 8316
rect 7466 8304 7472 8316
rect 7524 8304 7530 8356
rect 103330 7624 103336 7676
rect 103388 7664 103394 7676
rect 297358 7664 297364 7676
rect 103388 7636 297364 7664
rect 103388 7624 103394 7636
rect 297358 7624 297364 7636
rect 297416 7624 297422 7676
rect 47854 7556 47860 7608
rect 47912 7596 47918 7608
rect 275278 7596 275284 7608
rect 47912 7568 275284 7596
rect 47912 7556 47918 7568
rect 275278 7556 275284 7568
rect 275336 7556 275342 7608
rect 27706 6128 27712 6180
rect 27764 6168 27770 6180
rect 284938 6168 284944 6180
rect 27764 6140 284944 6168
rect 27764 6128 27770 6140
rect 284938 6128 284944 6140
rect 284996 6128 285002 6180
rect 56042 4768 56048 4820
rect 56100 4808 56106 4820
rect 268378 4808 268384 4820
rect 56100 4780 268384 4808
rect 56100 4768 56106 4780
rect 268378 4768 268384 4780
rect 268436 4768 268442 4820
rect 125870 3680 125876 3732
rect 125928 3720 125934 3732
rect 164878 3720 164884 3732
rect 125928 3692 164884 3720
rect 125928 3680 125934 3692
rect 164878 3680 164884 3692
rect 164936 3680 164942 3732
rect 110506 3612 110512 3664
rect 110564 3652 110570 3664
rect 110564 3624 111840 3652
rect 110564 3612 110570 3624
rect 67910 3544 67916 3596
rect 67968 3584 67974 3596
rect 67968 3556 74534 3584
rect 67968 3544 67974 3556
rect 2774 3476 2780 3528
rect 2832 3516 2838 3528
rect 3694 3516 3700 3528
rect 2832 3488 3700 3516
rect 2832 3476 2838 3488
rect 3694 3476 3700 3488
rect 3752 3476 3758 3528
rect 11054 3476 11060 3528
rect 11112 3516 11118 3528
rect 11974 3516 11980 3528
rect 11112 3488 11980 3516
rect 11112 3476 11118 3488
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 35894 3476 35900 3528
rect 35952 3516 35958 3528
rect 36814 3516 36820 3528
rect 35952 3488 36820 3516
rect 35952 3476 35958 3488
rect 36814 3476 36820 3488
rect 36872 3476 36878 3528
rect 44174 3476 44180 3528
rect 44232 3516 44238 3528
rect 45094 3516 45100 3528
rect 44232 3488 45100 3516
rect 44232 3476 44238 3488
rect 45094 3476 45100 3488
rect 45152 3476 45158 3528
rect 52454 3476 52460 3528
rect 52512 3516 52518 3528
rect 53374 3516 53380 3528
rect 52512 3488 53380 3516
rect 52512 3476 52518 3488
rect 53374 3476 53380 3488
rect 53432 3476 53438 3528
rect 69014 3476 69020 3528
rect 69072 3516 69078 3528
rect 69934 3516 69940 3528
rect 69072 3488 69940 3516
rect 69072 3476 69078 3488
rect 69934 3476 69940 3488
rect 69992 3476 69998 3528
rect 74506 3516 74534 3556
rect 110414 3544 110420 3596
rect 110472 3584 110478 3596
rect 111610 3584 111616 3596
rect 110472 3556 111616 3584
rect 110472 3544 110478 3556
rect 111610 3544 111616 3556
rect 111668 3544 111674 3596
rect 111812 3584 111840 3624
rect 112806 3612 112812 3664
rect 112864 3652 112870 3664
rect 206278 3652 206284 3664
rect 112864 3624 206284 3652
rect 112864 3612 112870 3624
rect 206278 3612 206284 3624
rect 206336 3612 206342 3664
rect 215938 3584 215944 3596
rect 111812 3556 215944 3584
rect 215938 3544 215944 3556
rect 215996 3544 216002 3596
rect 177298 3516 177304 3528
rect 74506 3488 177304 3516
rect 177298 3476 177304 3488
rect 177356 3476 177362 3528
rect 235810 3476 235816 3528
rect 235868 3516 235874 3528
rect 238018 3516 238024 3528
rect 235868 3488 238024 3516
rect 235868 3476 235874 3488
rect 238018 3476 238024 3488
rect 238076 3476 238082 3528
rect 23014 3408 23020 3460
rect 23072 3448 23078 3460
rect 47578 3448 47584 3460
rect 23072 3420 47584 3448
rect 23072 3408 23078 3420
rect 47578 3408 47584 3420
rect 47636 3408 47642 3460
rect 63218 3408 63224 3460
rect 63276 3448 63282 3460
rect 260098 3448 260104 3460
rect 63276 3420 260104 3448
rect 63276 3408 63282 3420
rect 260098 3408 260104 3420
rect 260156 3408 260162 3460
rect 118694 3340 118700 3392
rect 118752 3380 118758 3392
rect 119890 3380 119896 3392
rect 118752 3352 119896 3380
rect 118752 3340 118758 3352
rect 119890 3340 119896 3352
rect 119948 3340 119954 3392
rect 114002 2116 114008 2168
rect 114060 2156 114066 2168
rect 280798 2156 280804 2168
rect 114060 2128 280804 2156
rect 114060 2116 114066 2128
rect 280798 2116 280804 2128
rect 280856 2116 280862 2168
rect 109310 2048 109316 2100
rect 109368 2088 109374 2100
rect 295978 2088 295984 2100
rect 109368 2060 295984 2088
rect 109368 2048 109374 2060
rect 295978 2048 295984 2060
rect 296036 2048 296042 2100
<< via1 >>
rect 201500 703060 201552 703112
rect 202788 703060 202840 703112
rect 305644 703060 305696 703112
rect 494796 703060 494848 703112
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 87604 702992 87656 703044
rect 348792 702992 348844 703044
rect 107660 702924 107712 702976
rect 413652 702924 413704 702976
rect 129004 702856 129056 702908
rect 462320 702856 462372 702908
rect 53748 702788 53800 702840
rect 397460 702788 397512 702840
rect 106280 702720 106332 702772
rect 478512 702720 478564 702772
rect 57888 702652 57940 702704
rect 429844 702652 429896 702704
rect 124864 702584 124916 702636
rect 527180 702584 527232 702636
rect 133144 702516 133196 702568
rect 559656 702516 559708 702568
rect 79324 702448 79376 702500
rect 580908 702448 580960 702500
rect 55128 700340 55180 700392
rect 105452 700340 105504 700392
rect 75184 700272 75236 700324
rect 154120 700272 154172 700324
rect 24308 699660 24360 699712
rect 25504 699660 25556 699712
rect 214564 699660 214616 699712
rect 218980 699660 219032 699712
rect 359464 699660 359516 699712
rect 364984 699660 365036 699712
rect 151084 698912 151136 698964
rect 235172 698912 235224 698964
rect 62028 697620 62080 697672
rect 137836 697620 137888 697672
rect 266360 697620 266412 697672
rect 267648 697620 267700 697672
rect 134524 697552 134576 697604
rect 283840 697552 283892 697604
rect 126244 683136 126296 683188
rect 580172 683136 580224 683188
rect 3516 670692 3568 670744
rect 32404 670692 32456 670744
rect 148324 670692 148376 670744
rect 580172 670692 580224 670744
rect 3516 656888 3568 656940
rect 15844 656888 15896 656940
rect 123484 643084 123536 643136
rect 580172 643084 580224 643136
rect 3516 632068 3568 632120
rect 21364 632068 21416 632120
rect 3516 618264 3568 618316
rect 17224 618264 17276 618316
rect 130384 616836 130436 616888
rect 580172 616836 580224 616888
rect 3516 605820 3568 605872
rect 14464 605820 14516 605872
rect 52368 590656 52420 590708
rect 579804 590656 579856 590708
rect 3332 579640 3384 579692
rect 116584 579640 116636 579692
rect 142804 576852 142856 576904
rect 580172 576852 580224 576904
rect 3240 565836 3292 565888
rect 29644 565836 29696 565888
rect 97264 563048 97316 563100
rect 579804 563048 579856 563100
rect 3332 553392 3384 553444
rect 18604 553392 18656 553444
rect 123576 536800 123628 536852
rect 580172 536800 580224 536852
rect 2964 527144 3016 527196
rect 39304 527144 39356 527196
rect 141424 524424 141476 524476
rect 580172 524424 580224 524476
rect 66168 510620 66220 510672
rect 580172 510620 580224 510672
rect 3332 500964 3384 501016
rect 120080 500964 120132 501016
rect 126336 484372 126388 484424
rect 580172 484372 580224 484424
rect 3056 474716 3108 474768
rect 111064 474716 111116 474768
rect 124956 470568 125008 470620
rect 579988 470568 580040 470620
rect 3332 462340 3384 462392
rect 47584 462340 47636 462392
rect 3332 448536 3384 448588
rect 22744 448536 22796 448588
rect 129096 430584 129148 430636
rect 580172 430584 580224 430636
rect 2780 423512 2832 423564
rect 4804 423512 4856 423564
rect 93124 418140 93176 418192
rect 580172 418140 580224 418192
rect 3332 409844 3384 409896
rect 33784 409844 33836 409896
rect 67548 404336 67600 404388
rect 580172 404336 580224 404388
rect 3332 397468 3384 397520
rect 35164 397468 35216 397520
rect 127624 378156 127676 378208
rect 580172 378156 580224 378208
rect 3332 371220 3384 371272
rect 43444 371220 43496 371272
rect 3332 357416 3384 357468
rect 54484 357416 54536 357468
rect 76564 351908 76616 351960
rect 580172 351908 580224 351960
rect 3332 345040 3384 345092
rect 101404 345040 101456 345092
rect 88340 327700 88392 327752
rect 103796 327700 103848 327752
rect 3424 324912 3476 324964
rect 120264 324912 120316 324964
rect 91100 319404 91152 319456
rect 148324 319404 148376 319456
rect 3332 318792 3384 318844
rect 11704 318792 11756 318844
rect 116584 318724 116636 318776
rect 121460 318724 121512 318776
rect 11704 318044 11756 318096
rect 115940 318044 115992 318096
rect 93952 317500 94004 317552
rect 97264 317500 97316 317552
rect 3516 315256 3568 315308
rect 120172 315256 120224 315308
rect 77300 313896 77352 313948
rect 93124 313896 93176 313948
rect 54484 312536 54536 312588
rect 98000 312536 98052 312588
rect 125048 312536 125100 312588
rect 580264 312536 580316 312588
rect 14464 311108 14516 311160
rect 94136 311108 94188 311160
rect 101404 311108 101456 311160
rect 118700 311108 118752 311160
rect 15844 309748 15896 309800
rect 121552 309748 121604 309800
rect 123668 309748 123720 309800
rect 580172 309748 580224 309800
rect 71780 308388 71832 308440
rect 114560 308388 114612 308440
rect 122104 308388 122156 308440
rect 201500 308388 201552 308440
rect 63408 307776 63460 307828
rect 286324 307776 286376 307828
rect 89720 306348 89772 306400
rect 302884 306348 302936 306400
rect 69020 305600 69072 305652
rect 169760 305600 169812 305652
rect 92664 305056 92716 305108
rect 233884 305056 233936 305108
rect 3240 304988 3292 305040
rect 70400 304988 70452 305040
rect 75920 304988 75972 305040
rect 287704 304988 287756 305040
rect 25504 304240 25556 304292
rect 84476 304240 84528 304292
rect 85580 303764 85632 303816
rect 170404 303764 170456 303816
rect 81900 303696 81952 303748
rect 244924 303696 244976 303748
rect 74540 303628 74592 303680
rect 267740 303628 267792 303680
rect 90364 302404 90416 302456
rect 213184 302404 213236 302456
rect 69664 302336 69716 302388
rect 224224 302336 224276 302388
rect 100852 302268 100904 302320
rect 281540 302268 281592 302320
rect 71780 302200 71832 302252
rect 334624 302200 334676 302252
rect 22744 301452 22796 301504
rect 70400 301452 70452 301504
rect 121644 301452 121696 301504
rect 70400 301316 70452 301368
rect 85672 300908 85724 300960
rect 220084 300908 220136 300960
rect 102140 300840 102192 300892
rect 280160 300840 280212 300892
rect 102324 299684 102376 299736
rect 206284 299684 206336 299736
rect 84292 299616 84344 299668
rect 202144 299616 202196 299668
rect 70492 299548 70544 299600
rect 325792 299548 325844 299600
rect 80060 299480 80112 299532
rect 583024 299480 583076 299532
rect 4804 298732 4856 298784
rect 72608 298732 72660 298784
rect 89352 298460 89404 298512
rect 148324 298460 148376 298512
rect 110604 298392 110656 298444
rect 186964 298392 187016 298444
rect 79692 298324 79744 298376
rect 198004 298324 198056 298376
rect 83556 298256 83608 298308
rect 226984 298256 227036 298308
rect 111248 298188 111300 298240
rect 345112 298188 345164 298240
rect 73896 298120 73948 298172
rect 76564 298120 76616 298172
rect 88708 298120 88760 298172
rect 335360 298120 335412 298172
rect 112536 297032 112588 297084
rect 169024 297032 169076 297084
rect 82912 296964 82964 297016
rect 215944 296964 215996 297016
rect 117688 296896 117740 296948
rect 308404 296896 308456 296948
rect 113824 296828 113876 296880
rect 346400 296828 346452 296880
rect 97724 296760 97776 296812
rect 338120 296760 338172 296812
rect 77116 296692 77168 296744
rect 342904 296692 342956 296744
rect 99656 295672 99708 295724
rect 146944 295672 146996 295724
rect 11704 295604 11756 295656
rect 118332 295604 118384 295656
rect 88064 295536 88116 295588
rect 204904 295536 204956 295588
rect 68744 295468 68796 295520
rect 252560 295468 252612 295520
rect 75184 295400 75236 295452
rect 277400 295400 277452 295452
rect 99012 295332 99064 295384
rect 336740 295332 336792 295384
rect 85488 295060 85540 295112
rect 87604 295060 87656 295112
rect 73252 294584 73304 294636
rect 111800 294584 111852 294636
rect 70400 294312 70452 294364
rect 71044 294312 71096 294364
rect 77760 294312 77812 294364
rect 79324 294312 79376 294364
rect 85580 294312 85632 294364
rect 86500 294312 86552 294364
rect 93952 294312 94004 294364
rect 94780 294312 94832 294364
rect 106740 294312 106792 294364
rect 119712 294312 119764 294364
rect 67456 294244 67508 294296
rect 92572 294244 92624 294296
rect 111892 294244 111944 294296
rect 152464 294244 152516 294296
rect 87420 294176 87472 294228
rect 137284 294176 137336 294228
rect 91928 294108 91980 294160
rect 255412 294108 255464 294160
rect 3424 294040 3476 294092
rect 97080 294040 97132 294092
rect 114468 294040 114520 294092
rect 307024 294040 307076 294092
rect 50344 293972 50396 294024
rect 79048 293972 79100 294024
rect 81624 293972 81676 294024
rect 342260 293972 342312 294024
rect 111064 293224 111116 293276
rect 125600 293224 125652 293276
rect 2780 292816 2832 292868
rect 4804 292816 4856 292868
rect 8208 292816 8260 292868
rect 96436 292816 96488 292868
rect 109316 292816 109368 292868
rect 162124 292816 162176 292868
rect 53104 292748 53156 292800
rect 101588 292748 101640 292800
rect 103520 292748 103572 292800
rect 160744 292748 160796 292800
rect 93860 292680 93912 292732
rect 178684 292680 178736 292732
rect 80980 292612 81032 292664
rect 270500 292612 270552 292664
rect 68928 292544 68980 292596
rect 267832 292544 267884 292596
rect 119068 291932 119120 291984
rect 119804 291932 119856 291984
rect 115848 291864 115900 291916
rect 117228 291864 117280 291916
rect 3516 291796 3568 291848
rect 67456 291796 67508 291848
rect 155224 291320 155276 291372
rect 340880 291252 340932 291304
rect 69756 291184 69808 291236
rect 582748 291184 582800 291236
rect 121552 289892 121604 289944
rect 255320 289892 255372 289944
rect 25504 289824 25556 289876
rect 67640 289824 67692 289876
rect 121736 289824 121788 289876
rect 269120 289824 269172 289876
rect 121552 289756 121604 289808
rect 127624 289756 127676 289808
rect 121552 287036 121604 287088
rect 351920 287036 351972 287088
rect 32404 286968 32456 287020
rect 67640 286968 67692 287020
rect 122012 286288 122064 286340
rect 329840 286288 329892 286340
rect 59084 285676 59136 285728
rect 67732 285676 67784 285728
rect 63408 285608 63460 285660
rect 67640 285608 67692 285660
rect 121644 285540 121696 285592
rect 124956 285540 125008 285592
rect 121552 284316 121604 284368
rect 250444 284316 250496 284368
rect 121644 284180 121696 284232
rect 124864 284180 124916 284232
rect 57796 282888 57848 282940
rect 67640 282888 67692 282940
rect 121460 282888 121512 282940
rect 345020 282888 345072 282940
rect 121460 281596 121512 281648
rect 195244 281596 195296 281648
rect 121644 281528 121696 281580
rect 242164 281528 242216 281580
rect 121460 280236 121512 280288
rect 262220 280236 262272 280288
rect 63408 280168 63460 280220
rect 67640 280168 67692 280220
rect 121644 280168 121696 280220
rect 321560 280168 321612 280220
rect 66168 280100 66220 280152
rect 67732 280100 67784 280152
rect 121460 278808 121512 278860
rect 231124 278808 231176 278860
rect 51724 278740 51776 278792
rect 67640 278740 67692 278792
rect 121644 278740 121696 278792
rect 313924 278740 313976 278792
rect 56416 277448 56468 277500
rect 67640 277448 67692 277500
rect 121644 277448 121696 277500
rect 328460 277448 328512 277500
rect 54944 277380 54996 277432
rect 67732 277380 67784 277432
rect 121460 277380 121512 277432
rect 346492 277380 346544 277432
rect 65892 276088 65944 276140
rect 68008 276088 68060 276140
rect 55036 276020 55088 276072
rect 67640 276020 67692 276072
rect 121460 276020 121512 276072
rect 144184 276020 144236 276072
rect 122288 275272 122340 275324
rect 393964 275272 394016 275324
rect 57704 274660 57756 274712
rect 67640 274660 67692 274712
rect 121460 274660 121512 274712
rect 255504 274660 255556 274712
rect 17224 274592 17276 274644
rect 67732 274592 67784 274644
rect 121460 274252 121512 274304
rect 123668 274252 123720 274304
rect 66076 273232 66128 273284
rect 68008 273232 68060 273284
rect 121460 273232 121512 273284
rect 228364 273232 228416 273284
rect 61936 271940 61988 271992
rect 67640 271940 67692 271992
rect 60556 271872 60608 271924
rect 67732 271872 67784 271924
rect 130476 271872 130528 271924
rect 580172 271872 580224 271924
rect 121644 271124 121696 271176
rect 329932 271124 329984 271176
rect 49608 270512 49660 270564
rect 67640 270512 67692 270564
rect 6920 269764 6972 269816
rect 63500 269764 63552 269816
rect 59176 269084 59228 269136
rect 67640 269084 67692 269136
rect 121460 269084 121512 269136
rect 180064 269084 180116 269136
rect 121552 268336 121604 268388
rect 252652 268336 252704 268388
rect 32404 267724 32456 267776
rect 67640 267724 67692 267776
rect 121460 267724 121512 267776
rect 284944 267724 284996 267776
rect 29644 267656 29696 267708
rect 67732 267656 67784 267708
rect 63500 267588 63552 267640
rect 67640 267588 67692 267640
rect 121644 266976 121696 267028
rect 126336 266976 126388 267028
rect 121460 266432 121512 266484
rect 276664 266432 276716 266484
rect 121552 266364 121604 266416
rect 343732 266364 343784 266416
rect 21364 266296 21416 266348
rect 67732 266296 67784 266348
rect 121460 265004 121512 265056
rect 309784 265004 309836 265056
rect 53656 264936 53708 264988
rect 67640 264936 67692 264988
rect 121552 264936 121604 264988
rect 339592 264936 339644 264988
rect 59268 263644 59320 263696
rect 67640 263644 67692 263696
rect 17224 263576 17276 263628
rect 67732 263576 67784 263628
rect 121552 263576 121604 263628
rect 253940 263576 253992 263628
rect 18604 263508 18656 263560
rect 67640 263508 67692 263560
rect 121460 263508 121512 263560
rect 125600 263508 125652 263560
rect 144184 262828 144236 262880
rect 580356 262828 580408 262880
rect 60464 262216 60516 262268
rect 67640 262216 67692 262268
rect 121460 262216 121512 262268
rect 340880 262216 340932 262268
rect 119804 261468 119856 261520
rect 324596 261468 324648 261520
rect 65984 260924 66036 260976
rect 67640 260924 67692 260976
rect 61844 260856 61896 260908
rect 67732 260856 67784 260908
rect 121460 260856 121512 260908
rect 343640 260856 343692 260908
rect 39304 260788 39356 260840
rect 67640 260788 67692 260840
rect 56508 259428 56560 259480
rect 67640 259428 67692 259480
rect 121460 259428 121512 259480
rect 246304 259428 246356 259480
rect 121552 259360 121604 259412
rect 151084 259360 151136 259412
rect 342904 259360 342956 259412
rect 579804 259360 579856 259412
rect 64788 258136 64840 258188
rect 67640 258136 67692 258188
rect 57520 258068 57572 258120
rect 67732 258068 67784 258120
rect 121460 258068 121512 258120
rect 331220 258068 331272 258120
rect 121460 257864 121512 257916
rect 125048 257864 125100 257916
rect 50988 257320 51040 257372
rect 68284 257320 68336 257372
rect 124864 257320 124916 257372
rect 582380 257320 582432 257372
rect 14464 256708 14516 256760
rect 67640 256708 67692 256760
rect 121552 256708 121604 256760
rect 232504 256708 232556 256760
rect 121644 256640 121696 256692
rect 130384 256640 130436 256692
rect 121460 256572 121512 256624
rect 129096 256572 129148 256624
rect 64604 255348 64656 255400
rect 67640 255348 67692 255400
rect 60648 255280 60700 255332
rect 67732 255280 67784 255332
rect 57888 255212 57940 255264
rect 67640 255212 67692 255264
rect 121460 253988 121512 254040
rect 273260 253988 273312 254040
rect 3148 253920 3200 253972
rect 18604 253920 18656 253972
rect 121552 253920 121604 253972
rect 327080 253920 327132 253972
rect 64696 252628 64748 252680
rect 67640 252628 67692 252680
rect 22744 252560 22796 252612
rect 67732 252560 67784 252612
rect 121552 252560 121604 252612
rect 316684 252560 316736 252612
rect 121460 252492 121512 252544
rect 126244 252492 126296 252544
rect 63316 251200 63368 251252
rect 67640 251200 67692 251252
rect 121460 250452 121512 250504
rect 327172 250452 327224 250504
rect 60372 249840 60424 249892
rect 67640 249840 67692 249892
rect 58992 249772 59044 249824
rect 67732 249772 67784 249824
rect 121552 249772 121604 249824
rect 209044 249772 209096 249824
rect 62028 249704 62080 249756
rect 67640 249704 67692 249756
rect 121460 249704 121512 249756
rect 141424 249704 141476 249756
rect 67548 249636 67600 249688
rect 68376 249636 68428 249688
rect 57612 248412 57664 248464
rect 67640 248412 67692 248464
rect 121460 248412 121512 248464
rect 353300 248412 353352 248464
rect 62028 247120 62080 247172
rect 67640 247120 67692 247172
rect 61752 247052 61804 247104
rect 67732 247052 67784 247104
rect 121460 247052 121512 247104
rect 263600 247052 263652 247104
rect 53748 246984 53800 247036
rect 67640 246984 67692 247036
rect 64512 245624 64564 245676
rect 67732 245624 67784 245676
rect 121552 245624 121604 245676
rect 266452 245624 266504 245676
rect 33784 245556 33836 245608
rect 67640 245556 67692 245608
rect 121460 245556 121512 245608
rect 129004 245556 129056 245608
rect 121552 244332 121604 244384
rect 289084 244332 289136 244384
rect 63224 244264 63276 244316
rect 67640 244264 67692 244316
rect 128360 244264 128412 244316
rect 579896 244264 579948 244316
rect 4804 244196 4856 244248
rect 67732 244196 67784 244248
rect 121460 244196 121512 244248
rect 134524 244196 134576 244248
rect 122104 243516 122156 243568
rect 238024 243516 238076 243568
rect 121552 242836 121604 242888
rect 133144 242836 133196 242888
rect 121460 242768 121512 242820
rect 128360 242768 128412 242820
rect 160744 242224 160796 242276
rect 318064 242224 318116 242276
rect 121644 242156 121696 242208
rect 327264 242156 327316 242208
rect 63132 241476 63184 241528
rect 67640 241476 67692 241528
rect 121460 240184 121512 240236
rect 222844 240184 222896 240236
rect 3056 240116 3108 240168
rect 15200 240116 15252 240168
rect 121552 240116 121604 240168
rect 330024 240116 330076 240168
rect 118332 239912 118384 239964
rect 123484 239912 123536 239964
rect 73160 239776 73212 239828
rect 73884 239776 73936 239828
rect 75920 239776 75972 239828
rect 77104 239776 77156 239828
rect 77300 239776 77352 239828
rect 78392 239776 78444 239828
rect 78680 239776 78732 239828
rect 79680 239776 79732 239828
rect 82820 239776 82872 239828
rect 83544 239776 83596 239828
rect 86960 239776 87012 239828
rect 88052 239776 88104 239828
rect 89720 239776 89772 239828
rect 90628 239776 90680 239828
rect 92480 239776 92532 239828
rect 93204 239776 93256 239828
rect 104900 239776 104952 239828
rect 106084 239776 106136 239828
rect 114560 239776 114612 239828
rect 115744 239776 115796 239828
rect 64696 239504 64748 239556
rect 72424 239504 72476 239556
rect 63316 239436 63368 239488
rect 98644 239436 98696 239488
rect 3608 239368 3660 239420
rect 63500 239368 63552 239420
rect 69664 239368 69716 239420
rect 312544 239368 312596 239420
rect 84292 239300 84344 239352
rect 85488 239300 85540 239352
rect 106740 238756 106792 238808
rect 266360 238756 266412 238808
rect 15200 238688 15252 238740
rect 103520 238688 103572 238740
rect 113824 238688 113876 238740
rect 305644 238688 305696 238740
rect 40040 238620 40092 238672
rect 95792 238620 95844 238672
rect 117044 238620 117096 238672
rect 124864 238620 124916 238672
rect 52368 238552 52420 238604
rect 75828 238552 75880 238604
rect 91284 238552 91336 238604
rect 130476 238552 130528 238604
rect 63500 238484 63552 238536
rect 86776 238484 86828 238536
rect 115112 238484 115164 238536
rect 123576 238484 123628 238536
rect 102876 238212 102928 238264
rect 106924 238212 106976 238264
rect 81624 238144 81676 238196
rect 114836 238144 114888 238196
rect 72608 238076 72660 238128
rect 91100 238076 91152 238128
rect 105452 238076 105504 238128
rect 196624 238076 196676 238128
rect 71320 238008 71372 238060
rect 79324 238008 79376 238060
rect 86132 238008 86184 238060
rect 582380 238008 582432 238060
rect 35164 237328 35216 237380
rect 82268 237328 82320 237380
rect 98368 237328 98420 237380
rect 359464 237328 359516 237380
rect 47584 237260 47636 237312
rect 114468 237260 114520 237312
rect 55128 237192 55180 237244
rect 89352 237192 89404 237244
rect 67364 236648 67416 236700
rect 214656 236648 214708 236700
rect 18604 235900 18656 235952
rect 112536 235900 112588 235952
rect 43444 235832 43496 235884
rect 99012 235832 99064 235884
rect 80336 235288 80388 235340
rect 320824 235288 320876 235340
rect 117688 235220 117740 235272
rect 583116 235220 583168 235272
rect 91928 234540 91980 234592
rect 582656 234540 582708 234592
rect 69020 233928 69072 233980
rect 69756 233928 69808 233980
rect 63224 233860 63276 233912
rect 191196 233860 191248 233912
rect 93860 233724 93912 233776
rect 94044 233724 94096 233776
rect 114836 233180 114888 233232
rect 214564 233180 214616 233232
rect 69204 232500 69256 232552
rect 251180 232500 251232 232552
rect 84108 231820 84160 231872
rect 84844 231820 84896 231872
rect 106832 231752 106884 231804
rect 542360 231752 542412 231804
rect 60372 231208 60424 231260
rect 160744 231208 160796 231260
rect 15844 231140 15896 231192
rect 109868 231140 109920 231192
rect 111800 231140 111852 231192
rect 276020 231140 276072 231192
rect 108580 231072 108632 231124
rect 328552 231072 328604 231124
rect 91100 230392 91152 230444
rect 582564 230392 582616 230444
rect 67272 228420 67324 228472
rect 315304 228420 315356 228472
rect 76012 228352 76064 228404
rect 582564 228352 582616 228404
rect 54944 225564 54996 225616
rect 305644 225564 305696 225616
rect 82912 224272 82964 224324
rect 184204 224272 184256 224324
rect 97632 224204 97684 224256
rect 342352 224204 342404 224256
rect 84292 222844 84344 222896
rect 254124 222844 254176 222896
rect 89812 221484 89864 221536
rect 252744 221484 252796 221536
rect 61844 221416 61896 221468
rect 334072 221416 334124 221468
rect 1308 220192 1360 220244
rect 119804 220192 119856 220244
rect 115940 220124 115992 220176
rect 259736 220124 259788 220176
rect 113364 220056 113416 220108
rect 304264 220056 304316 220108
rect 77392 218696 77444 218748
rect 330116 218696 330168 218748
rect 137284 217404 137336 217456
rect 245016 217404 245068 217456
rect 53656 217336 53708 217388
rect 298744 217336 298796 217388
rect 75920 217268 75972 217320
rect 321652 217268 321704 217320
rect 78772 215976 78824 216028
rect 273352 215976 273404 216028
rect 94044 215908 94096 215960
rect 300124 215908 300176 215960
rect 3332 215228 3384 215280
rect 17224 215228 17276 215280
rect 100852 214616 100904 214668
rect 254032 214616 254084 214668
rect 74632 214548 74684 214600
rect 323124 214548 323176 214600
rect 60464 213188 60516 213240
rect 233976 213188 234028 213240
rect 110512 211828 110564 211880
rect 238116 211828 238168 211880
rect 96620 211760 96672 211812
rect 260932 211760 260984 211812
rect 146944 210468 146996 210520
rect 271880 210468 271932 210520
rect 61752 210400 61804 210452
rect 240784 210400 240836 210452
rect 93952 209108 94004 209160
rect 278780 209108 278832 209160
rect 61936 209040 61988 209092
rect 270684 209040 270736 209092
rect 56416 207748 56468 207800
rect 264980 207748 265032 207800
rect 57612 207680 57664 207732
rect 277492 207680 277544 207732
rect 78680 207612 78732 207664
rect 335452 207612 335504 207664
rect 127716 206932 127768 206984
rect 580172 206932 580224 206984
rect 77300 206320 77352 206372
rect 263692 206320 263744 206372
rect 98644 206252 98696 206304
rect 332876 206252 332928 206304
rect 103612 205028 103664 205080
rect 191104 205028 191156 205080
rect 148324 204960 148376 205012
rect 343824 204960 343876 205012
rect 63408 204892 63460 204944
rect 266360 204892 266412 204944
rect 100760 203600 100812 203652
rect 261116 203600 261168 203652
rect 155224 203532 155276 203584
rect 339776 203532 339828 203584
rect 3056 202784 3108 202836
rect 120080 202784 120132 202836
rect 103704 202172 103756 202224
rect 216036 202172 216088 202224
rect 104900 202104 104952 202156
rect 340972 202104 341024 202156
rect 59176 200744 59228 200796
rect 271972 200744 272024 200796
rect 250444 199588 250496 199640
rect 338396 199588 338448 199640
rect 57704 199520 57756 199572
rect 258080 199520 258132 199572
rect 60556 199452 60608 199504
rect 276112 199452 276164 199504
rect 87052 199384 87104 199436
rect 323032 199384 323084 199436
rect 89720 198024 89772 198076
rect 254216 198024 254268 198076
rect 63132 197956 63184 198008
rect 262312 197956 262364 198008
rect 99472 196596 99524 196648
rect 249800 196596 249852 196648
rect 86960 195304 87012 195356
rect 267924 195304 267976 195356
rect 99380 195236 99432 195288
rect 328644 195236 328696 195288
rect 66076 194080 66128 194132
rect 251272 194080 251324 194132
rect 57520 194012 57572 194064
rect 273444 194012 273496 194064
rect 65984 193944 66036 193996
rect 324412 193944 324464 193996
rect 88432 193876 88484 193928
rect 347872 193876 347924 193928
rect 64512 193808 64564 193860
rect 347964 193808 348016 193860
rect 574744 193128 574796 193180
rect 580172 193128 580224 193180
rect 106924 192448 106976 192500
rect 259552 192448 259604 192500
rect 92572 191360 92624 191412
rect 249892 191360 249944 191412
rect 84200 191292 84252 191344
rect 321744 191292 321796 191344
rect 107660 191224 107712 191276
rect 347780 191224 347832 191276
rect 95332 191156 95384 191208
rect 336832 191156 336884 191208
rect 102140 191088 102192 191140
rect 343916 191088 343968 191140
rect 169024 189796 169076 189848
rect 269212 189796 269264 189848
rect 73160 189728 73212 189780
rect 325884 189728 325936 189780
rect 106188 189048 106240 189100
rect 173164 189048 173216 189100
rect 160744 188572 160796 188624
rect 274732 188572 274784 188624
rect 214656 188504 214708 188556
rect 334164 188504 334216 188556
rect 55036 188436 55088 188488
rect 259644 188436 259696 188488
rect 64788 188368 64840 188420
rect 270592 188368 270644 188420
rect 70400 188300 70452 188352
rect 345204 188300 345256 188352
rect 107568 187756 107620 187808
rect 171784 187756 171836 187808
rect 133788 187688 133840 187740
rect 214564 187688 214616 187740
rect 206284 187008 206336 187060
rect 274640 187008 274692 187060
rect 17224 186940 17276 186992
rect 110420 186940 110472 186992
rect 152464 186940 152516 186992
rect 331312 186940 331364 186992
rect 132408 186464 132460 186516
rect 170588 186464 170640 186516
rect 100668 186396 100720 186448
rect 169024 186396 169076 186448
rect 118608 186328 118660 186380
rect 214656 186328 214708 186380
rect 118700 185852 118752 185904
rect 346584 185852 346636 185904
rect 80060 185784 80112 185836
rect 327356 185784 327408 185836
rect 65892 185716 65944 185768
rect 324504 185716 324556 185768
rect 67548 185648 67600 185700
rect 334256 185648 334308 185700
rect 58992 185580 59044 185632
rect 331404 185580 331456 185632
rect 121368 184900 121420 184952
rect 170496 184900 170548 184952
rect 180064 184288 180116 184340
rect 262404 184288 262456 184340
rect 289084 184288 289136 184340
rect 338212 184288 338264 184340
rect 57796 184220 57848 184272
rect 308496 184220 308548 184272
rect 69020 184152 69072 184204
rect 323216 184152 323268 184204
rect 114468 183540 114520 183592
rect 169300 183540 169352 183592
rect 244924 183132 244976 183184
rect 256792 183132 256844 183184
rect 238116 183064 238168 183116
rect 256976 183064 257028 183116
rect 213184 182996 213236 183048
rect 265072 182996 265124 183048
rect 186964 182928 187016 182980
rect 262496 182928 262548 182980
rect 276664 182928 276716 182980
rect 336924 182928 336976 182980
rect 93860 182860 93912 182912
rect 338488 182860 338540 182912
rect 56508 182792 56560 182844
rect 345296 182792 345348 182844
rect 116952 182316 117004 182368
rect 167736 182316 167788 182368
rect 97540 182248 97592 182300
rect 169208 182248 169260 182300
rect 129464 182180 129516 182232
rect 213276 182180 213328 182232
rect 316684 181636 316736 181688
rect 342536 181636 342588 181688
rect 202144 181568 202196 181620
rect 246948 181568 247000 181620
rect 300124 181568 300176 181620
rect 332692 181568 332744 181620
rect 170404 181500 170456 181552
rect 316316 181500 316368 181552
rect 318064 181500 318116 181552
rect 341156 181500 341208 181552
rect 74724 181432 74776 181484
rect 252836 181432 252888 181484
rect 307024 181432 307076 181484
rect 339684 181432 339736 181484
rect 112996 180820 113048 180872
rect 166356 180820 166408 180872
rect 238024 180412 238076 180464
rect 261024 180412 261076 180464
rect 228364 180344 228416 180396
rect 259460 180344 259512 180396
rect 222844 180276 222896 180328
rect 258172 180276 258224 180328
rect 191196 180208 191248 180260
rect 255596 180208 255648 180260
rect 72424 180140 72476 180192
rect 332784 180140 332836 180192
rect 67456 180072 67508 180124
rect 335544 180072 335596 180124
rect 123760 179460 123812 179512
rect 167828 179460 167880 179512
rect 128084 179392 128136 179444
rect 211804 179392 211856 179444
rect 287704 179324 287756 179376
rect 338304 179324 338356 179376
rect 231124 178916 231176 178968
rect 249064 178916 249116 178968
rect 209044 178848 209096 178900
rect 249248 178848 249300 178900
rect 215944 178780 215996 178832
rect 258264 178780 258316 178832
rect 204904 178712 204956 178764
rect 260840 178712 260892 178764
rect 162124 178644 162176 178696
rect 331496 178644 331548 178696
rect 148232 178304 148284 178356
rect 169116 178304 169168 178356
rect 134800 178236 134852 178288
rect 165344 178236 165396 178288
rect 126060 178168 126112 178220
rect 167920 178168 167972 178220
rect 115848 178100 115900 178152
rect 166448 178100 166500 178152
rect 109960 178032 110012 178084
rect 170404 178032 170456 178084
rect 242164 177964 242216 178016
rect 249156 177964 249208 178016
rect 312544 177488 312596 177540
rect 332600 177488 332652 177540
rect 246304 177420 246356 177472
rect 263784 177420 263836 177472
rect 315304 177420 315356 177472
rect 335636 177420 335688 177472
rect 233976 177352 234028 177404
rect 258356 177352 258408 177404
rect 304264 177352 304316 177404
rect 333980 177352 334032 177404
rect 4804 177284 4856 177336
rect 82820 177284 82872 177336
rect 195244 177284 195296 177336
rect 251364 177284 251416 177336
rect 284944 177284 284996 177336
rect 337016 177284 337068 177336
rect 130752 177012 130804 177064
rect 165528 177012 165580 177064
rect 104624 176944 104676 176996
rect 165436 176944 165488 176996
rect 103336 176876 103388 176928
rect 167644 176876 167696 176928
rect 136088 176808 136140 176860
rect 213920 176808 213972 176860
rect 124496 176740 124548 176792
rect 211896 176740 211948 176792
rect 108120 176672 108172 176724
rect 195336 176672 195388 176724
rect 305644 176604 305696 176656
rect 321468 176604 321520 176656
rect 158904 176264 158956 176316
rect 166264 176264 166316 176316
rect 121920 176196 121972 176248
rect 166540 176196 166592 176248
rect 113180 176128 113232 176180
rect 170680 176128 170732 176180
rect 128176 176060 128228 176112
rect 212264 176060 212316 176112
rect 119436 175992 119488 176044
rect 214748 175992 214800 176044
rect 240784 175992 240836 176044
rect 256700 175992 256752 176044
rect 338396 175992 338448 176044
rect 100760 175924 100812 175976
rect 209044 175924 209096 175976
rect 233884 175924 233936 175976
rect 249984 175924 250036 175976
rect 313924 175924 313976 175976
rect 321468 175924 321520 175976
rect 338396 175788 338448 175840
rect 165344 175176 165396 175228
rect 213920 175176 213972 175228
rect 165528 174496 165580 174548
rect 214012 174496 214064 174548
rect 287796 174020 287848 174072
rect 307576 174020 307628 174072
rect 268384 173952 268436 174004
rect 307668 173952 307720 174004
rect 264244 173884 264296 173936
rect 306564 173884 306616 173936
rect 170588 173816 170640 173868
rect 213920 173816 213972 173868
rect 165436 173136 165488 173188
rect 214656 173136 214708 173188
rect 284944 172660 284996 172712
rect 307484 172660 307536 172712
rect 276664 172592 276716 172644
rect 307576 172592 307628 172644
rect 252468 172524 252520 172576
rect 259644 172524 259696 172576
rect 267188 172524 267240 172576
rect 307668 172524 307720 172576
rect 212264 172456 212316 172508
rect 213920 172456 213972 172508
rect 324320 172456 324372 172508
rect 336832 172456 336884 172508
rect 252468 172320 252520 172372
rect 263600 172320 263652 172372
rect 252376 171368 252428 171420
rect 259460 171368 259512 171420
rect 289176 171232 289228 171284
rect 306564 171232 306616 171284
rect 265808 171164 265860 171216
rect 307576 171164 307628 171216
rect 168012 171096 168064 171148
rect 214472 171096 214524 171148
rect 260288 171096 260340 171148
rect 307668 171096 307720 171148
rect 167920 171028 167972 171080
rect 213920 171028 213972 171080
rect 324320 171028 324372 171080
rect 338120 171028 338172 171080
rect 211804 170960 211856 171012
rect 214472 170960 214524 171012
rect 252468 170756 252520 170808
rect 256700 170756 256752 170808
rect 286416 169872 286468 169924
rect 306564 169872 306616 169924
rect 252468 169804 252520 169856
rect 258080 169804 258132 169856
rect 265716 169804 265768 169856
rect 307576 169804 307628 169856
rect 259000 169736 259052 169788
rect 307668 169736 307720 169788
rect 167828 169668 167880 169720
rect 213920 169668 213972 169720
rect 252376 169668 252428 169720
rect 260932 169668 260984 169720
rect 211896 169600 211948 169652
rect 214012 169600 214064 169652
rect 252284 169600 252336 169652
rect 260840 169600 260892 169652
rect 252468 168920 252520 168972
rect 259552 168920 259604 168972
rect 291844 168512 291896 168564
rect 307668 168512 307720 168564
rect 269856 168444 269908 168496
rect 307484 168444 307536 168496
rect 261576 168376 261628 168428
rect 307576 168376 307628 168428
rect 166540 168308 166592 168360
rect 213920 168308 213972 168360
rect 252376 168308 252428 168360
rect 261024 168308 261076 168360
rect 324320 168308 324372 168360
rect 332784 168308 332836 168360
rect 170496 168240 170548 168292
rect 214012 168240 214064 168292
rect 252284 168240 252336 168292
rect 255412 168240 255464 168292
rect 324412 168240 324464 168292
rect 332600 168240 332652 168292
rect 252468 167832 252520 167884
rect 258264 167832 258316 167884
rect 282276 167152 282328 167204
rect 307668 167152 307720 167204
rect 271328 167084 271380 167136
rect 307576 167084 307628 167136
rect 261668 167016 261720 167068
rect 307484 167016 307536 167068
rect 167736 166948 167788 167000
rect 213920 166948 213972 167000
rect 324320 166948 324372 167000
rect 335636 166948 335688 167000
rect 252468 166200 252520 166252
rect 258172 166200 258224 166252
rect 252376 165724 252428 165776
rect 258356 165724 258408 165776
rect 280804 165724 280856 165776
rect 307668 165724 307720 165776
rect 272616 165656 272668 165708
rect 307300 165656 307352 165708
rect 258908 165588 258960 165640
rect 307576 165588 307628 165640
rect 166448 165520 166500 165572
rect 213920 165520 213972 165572
rect 252376 165520 252428 165572
rect 264980 165520 265032 165572
rect 324320 165520 324372 165572
rect 343916 165520 343968 165572
rect 169300 165452 169352 165504
rect 214012 165452 214064 165504
rect 252468 165452 252520 165504
rect 262496 165452 262548 165504
rect 300400 164364 300452 164416
rect 307576 164364 307628 164416
rect 274088 164296 274140 164348
rect 307668 164296 307720 164348
rect 258816 164228 258868 164280
rect 307300 164228 307352 164280
rect 3240 164160 3292 164212
rect 50344 164160 50396 164212
rect 166356 164160 166408 164212
rect 214012 164160 214064 164212
rect 252468 164160 252520 164212
rect 267740 164160 267792 164212
rect 324412 164160 324464 164212
rect 345296 164160 345348 164212
rect 170680 164092 170732 164144
rect 213920 164092 213972 164144
rect 251456 164092 251508 164144
rect 253940 164092 253992 164144
rect 324320 164092 324372 164144
rect 334072 164092 334124 164144
rect 297456 163004 297508 163056
rect 307576 163004 307628 163056
rect 269764 162936 269816 162988
rect 307484 162936 307536 162988
rect 261484 162868 261536 162920
rect 307668 162868 307720 162920
rect 170404 162800 170456 162852
rect 213920 162800 213972 162852
rect 252376 162800 252428 162852
rect 266360 162800 266412 162852
rect 324320 162800 324372 162852
rect 331496 162800 331548 162852
rect 252284 162732 252336 162784
rect 263692 162732 263744 162784
rect 252468 162664 252520 162716
rect 262404 162664 262456 162716
rect 324320 161848 324372 161900
rect 327264 161848 327316 161900
rect 289360 161576 289412 161628
rect 307576 161576 307628 161628
rect 286324 161508 286376 161560
rect 307668 161508 307720 161560
rect 253204 161440 253256 161492
rect 307484 161440 307536 161492
rect 171784 161372 171836 161424
rect 214012 161372 214064 161424
rect 324320 161372 324372 161424
rect 345112 161372 345164 161424
rect 195336 161304 195388 161356
rect 213920 161304 213972 161356
rect 324412 161304 324464 161356
rect 338396 161304 338448 161356
rect 252468 160760 252520 160812
rect 259736 160760 259788 160812
rect 267280 160692 267332 160744
rect 307300 160692 307352 160744
rect 304540 160148 304592 160200
rect 307668 160148 307720 160200
rect 260104 160080 260156 160132
rect 307576 160080 307628 160132
rect 173164 160012 173216 160064
rect 213920 160012 213972 160064
rect 252468 160012 252520 160064
rect 267832 160012 267884 160064
rect 324320 160012 324372 160064
rect 345204 160012 345256 160064
rect 252008 159944 252060 159996
rect 255320 159944 255372 159996
rect 298744 158856 298796 158908
rect 306564 158856 306616 158908
rect 262956 158788 263008 158840
rect 307300 158788 307352 158840
rect 258724 158720 258776 158772
rect 307668 158720 307720 158772
rect 167644 158652 167696 158704
rect 213920 158652 213972 158704
rect 324412 158652 324464 158704
rect 341156 158652 341208 158704
rect 186964 158584 187016 158636
rect 214012 158584 214064 158636
rect 324320 158584 324372 158636
rect 336924 158584 336976 158636
rect 256148 157564 256200 157616
rect 306932 157564 306984 157616
rect 295984 157496 296036 157548
rect 307668 157496 307720 157548
rect 267096 157428 267148 157480
rect 307576 157428 307628 157480
rect 169024 157292 169076 157344
rect 214012 157292 214064 157344
rect 252468 157292 252520 157344
rect 281540 157292 281592 157344
rect 324320 157292 324372 157344
rect 328644 157292 328696 157344
rect 209044 157224 209096 157276
rect 213920 157224 213972 157276
rect 252376 157224 252428 157276
rect 270684 157224 270736 157276
rect 252468 157156 252520 157208
rect 263784 157156 263836 157208
rect 296168 156068 296220 156120
rect 307668 156068 307720 156120
rect 262864 156000 262916 156052
rect 307484 156000 307536 156052
rect 260196 155932 260248 155984
rect 307576 155932 307628 155984
rect 169208 155864 169260 155916
rect 213920 155864 213972 155916
rect 252376 155864 252428 155916
rect 265072 155864 265124 155916
rect 324412 155864 324464 155916
rect 347964 155864 348016 155916
rect 252468 155796 252520 155848
rect 261116 155796 261168 155848
rect 324320 155796 324372 155848
rect 346492 155796 346544 155848
rect 251456 155728 251508 155780
rect 254124 155728 254176 155780
rect 300216 154708 300268 154760
rect 307668 154708 307720 154760
rect 285036 154640 285088 154692
rect 306564 154640 306616 154692
rect 264520 154572 264572 154624
rect 307300 154572 307352 154624
rect 252376 154504 252428 154556
rect 271972 154504 272024 154556
rect 324320 154504 324372 154556
rect 347872 154504 347924 154556
rect 252468 154436 252520 154488
rect 267924 154436 267976 154488
rect 252284 154368 252336 154420
rect 255504 154368 255556 154420
rect 324320 153756 324372 153808
rect 327356 153756 327408 153808
rect 198004 153280 198056 153332
rect 214012 153280 214064 153332
rect 303528 153280 303580 153332
rect 307668 153280 307720 153332
rect 178684 153212 178736 153264
rect 213920 153212 213972 153264
rect 282460 153212 282512 153264
rect 306564 153212 306616 153264
rect 324412 153144 324464 153196
rect 342536 153144 342588 153196
rect 393964 153144 394016 153196
rect 579804 153144 579856 153196
rect 252468 153076 252520 153128
rect 269212 153076 269264 153128
rect 304264 151920 304316 151972
rect 307576 151920 307628 151972
rect 268476 151852 268528 151904
rect 307668 151852 307720 151904
rect 177580 151784 177632 151836
rect 213920 151784 213972 151836
rect 256056 151784 256108 151836
rect 307484 151784 307536 151836
rect 252468 151716 252520 151768
rect 276020 151716 276072 151768
rect 324320 151648 324372 151700
rect 347780 151648 347832 151700
rect 252008 151444 252060 151496
rect 254216 151444 254268 151496
rect 173256 151036 173308 151088
rect 214380 151036 214432 151088
rect 287980 150560 288032 150612
rect 307668 150560 307720 150612
rect 264336 150492 264388 150544
rect 307300 150492 307352 150544
rect 175924 150424 175976 150476
rect 214012 150424 214064 150476
rect 254584 150424 254636 150476
rect 306932 150424 306984 150476
rect 3516 150356 3568 150408
rect 25504 150356 25556 150408
rect 169116 150356 169168 150408
rect 213920 150356 213972 150408
rect 252468 150356 252520 150408
rect 278780 150356 278832 150408
rect 324320 150356 324372 150408
rect 334256 150356 334308 150408
rect 252376 150288 252428 150340
rect 273260 150288 273312 150340
rect 252284 150220 252336 150272
rect 256792 150220 256844 150272
rect 324412 150220 324464 150272
rect 327172 150220 327224 150272
rect 299112 149744 299164 149796
rect 306656 149744 306708 149796
rect 257344 149676 257396 149728
rect 307116 149676 307168 149728
rect 281080 149064 281132 149116
rect 307668 149064 307720 149116
rect 166264 148996 166316 149048
rect 213920 148996 213972 149048
rect 252468 148996 252520 149048
rect 280160 148996 280212 149048
rect 324320 148996 324372 149048
rect 343732 148996 343784 149048
rect 252376 148928 252428 148980
rect 276112 148928 276164 148980
rect 264428 147772 264480 147824
rect 306564 147772 306616 147824
rect 167736 147636 167788 147688
rect 213920 147636 213972 147688
rect 301780 147636 301832 147688
rect 307668 147636 307720 147688
rect 252468 147568 252520 147620
rect 274732 147568 274784 147620
rect 324320 147568 324372 147620
rect 335360 147568 335412 147620
rect 251272 147500 251324 147552
rect 254032 147500 254084 147552
rect 290648 146888 290700 146940
rect 307208 146888 307260 146940
rect 210424 146344 210476 146396
rect 214012 146344 214064 146396
rect 255964 146344 256016 146396
rect 307300 146344 307352 146396
rect 174544 146276 174596 146328
rect 213920 146276 213972 146328
rect 254676 146276 254728 146328
rect 306932 146276 306984 146328
rect 252284 146208 252336 146260
rect 273352 146208 273404 146260
rect 324320 146208 324372 146260
rect 339776 146208 339828 146260
rect 252468 146140 252520 146192
rect 273444 146140 273496 146192
rect 324412 146140 324464 146192
rect 328736 146140 328788 146192
rect 252376 146072 252428 146124
rect 262312 146072 262364 146124
rect 292120 145596 292172 145648
rect 307576 145596 307628 145648
rect 252008 145528 252060 145580
rect 264244 145528 264296 145580
rect 285220 145528 285272 145580
rect 307484 145528 307536 145580
rect 173164 144984 173216 145036
rect 214012 144984 214064 145036
rect 169024 144916 169076 144968
rect 213920 144916 213972 144968
rect 252468 144848 252520 144900
rect 266452 144848 266504 144900
rect 324320 144848 324372 144900
rect 331404 144848 331456 144900
rect 324412 144780 324464 144832
rect 329932 144780 329984 144832
rect 299020 143692 299072 143744
rect 307484 143692 307536 143744
rect 202144 143624 202196 143676
rect 213920 143624 213972 143676
rect 268568 143624 268620 143676
rect 307576 143624 307628 143676
rect 166264 143556 166316 143608
rect 214012 143556 214064 143608
rect 253296 143556 253348 143608
rect 307668 143556 307720 143608
rect 252376 143488 252428 143540
rect 270500 143488 270552 143540
rect 324412 143488 324464 143540
rect 351920 143488 351972 143540
rect 252468 143420 252520 143472
rect 269120 143420 269172 143472
rect 324320 143420 324372 143472
rect 334164 143420 334216 143472
rect 251916 142808 251968 142860
rect 280804 142808 280856 142860
rect 300308 142264 300360 142316
rect 307668 142264 307720 142316
rect 280988 142196 281040 142248
rect 306564 142196 306616 142248
rect 206376 142128 206428 142180
rect 213920 142128 213972 142180
rect 269948 142128 270000 142180
rect 307576 142128 307628 142180
rect 252468 142060 252520 142112
rect 262220 142060 262272 142112
rect 324412 142060 324464 142112
rect 342260 142060 342312 142112
rect 324320 141992 324372 142044
rect 339592 141992 339644 142044
rect 253388 141380 253440 141432
rect 307484 141380 307536 141432
rect 275284 140904 275336 140956
rect 307668 140904 307720 140956
rect 177396 140836 177448 140888
rect 213920 140836 213972 140888
rect 294880 140836 294932 140888
rect 306564 140836 306616 140888
rect 167644 140768 167696 140820
rect 214012 140768 214064 140820
rect 304448 140768 304500 140820
rect 307576 140768 307628 140820
rect 252468 140700 252520 140752
rect 274640 140700 274692 140752
rect 324320 140700 324372 140752
rect 329840 140700 329892 140752
rect 252376 140632 252428 140684
rect 256976 140632 257028 140684
rect 257436 140020 257488 140072
rect 307116 140020 307168 140072
rect 209044 139476 209096 139528
rect 213920 139476 213972 139528
rect 289084 139476 289136 139528
rect 306932 139476 306984 139528
rect 171784 139408 171836 139460
rect 214012 139408 214064 139460
rect 279516 139408 279568 139460
rect 307300 139408 307352 139460
rect 252284 139340 252336 139392
rect 255596 139340 255648 139392
rect 324412 139340 324464 139392
rect 332876 139340 332928 139392
rect 324320 139272 324372 139324
rect 331312 139272 331364 139324
rect 252192 138660 252244 138712
rect 265808 138660 265860 138712
rect 280804 138116 280856 138168
rect 307668 138116 307720 138168
rect 267004 138048 267056 138100
rect 307576 138048 307628 138100
rect 170404 137980 170456 138032
rect 213920 137980 213972 138032
rect 250444 137980 250496 138032
rect 306564 137980 306616 138032
rect 3516 137912 3568 137964
rect 14464 137912 14516 137964
rect 252284 137912 252336 137964
rect 277492 137912 277544 137964
rect 324320 137912 324372 137964
rect 343640 137912 343692 137964
rect 252376 137844 252428 137896
rect 277400 137844 277452 137896
rect 324412 137844 324464 137896
rect 335452 137844 335504 137896
rect 252468 137776 252520 137828
rect 271880 137776 271932 137828
rect 251824 137300 251876 137352
rect 295984 137300 296036 137352
rect 171968 137232 172020 137284
rect 214564 137232 214616 137284
rect 253480 137232 253532 137284
rect 307024 137232 307076 137284
rect 297364 136688 297416 136740
rect 307668 136688 307720 136740
rect 204904 136620 204956 136672
rect 213920 136620 213972 136672
rect 293224 136620 293276 136672
rect 307576 136620 307628 136672
rect 252284 136552 252336 136604
rect 287796 136552 287848 136604
rect 324320 136552 324372 136604
rect 341064 136552 341116 136604
rect 252468 136484 252520 136536
rect 270592 136484 270644 136536
rect 252376 136416 252428 136468
rect 268384 136416 268436 136468
rect 324964 136212 325016 136264
rect 327080 136212 327132 136264
rect 302884 135464 302936 135516
rect 307300 135464 307352 135516
rect 287704 135396 287756 135448
rect 306564 135396 306616 135448
rect 195244 135328 195296 135380
rect 214012 135328 214064 135380
rect 283564 135328 283616 135380
rect 307484 135328 307536 135380
rect 170496 135260 170548 135312
rect 213920 135260 213972 135312
rect 278136 135260 278188 135312
rect 307668 135260 307720 135312
rect 252468 135192 252520 135244
rect 276664 135192 276716 135244
rect 307208 135192 307260 135244
rect 307484 135192 307536 135244
rect 252376 135124 252428 135176
rect 267188 135124 267240 135176
rect 324320 135124 324372 135176
rect 339500 135124 339552 135176
rect 177488 133968 177540 134020
rect 213920 133968 213972 134020
rect 291936 133968 291988 134020
rect 307576 133968 307628 134020
rect 167828 133900 167880 133952
rect 214012 133900 214064 133952
rect 276756 133900 276808 133952
rect 307668 133900 307720 133952
rect 252376 133832 252428 133884
rect 289176 133832 289228 133884
rect 324320 133832 324372 133884
rect 330024 133832 330076 133884
rect 252468 133764 252520 133816
rect 284944 133764 284996 133816
rect 286600 133152 286652 133204
rect 306748 133152 306800 133204
rect 196716 132540 196768 132592
rect 214012 132540 214064 132592
rect 290556 132540 290608 132592
rect 307668 132540 307720 132592
rect 173348 132472 173400 132524
rect 213920 132472 213972 132524
rect 282184 132472 282236 132524
rect 307576 132472 307628 132524
rect 252284 132404 252336 132456
rect 286416 132404 286468 132456
rect 324412 132404 324464 132456
rect 346400 132404 346452 132456
rect 252468 132336 252520 132388
rect 265716 132336 265768 132388
rect 324320 132336 324372 132388
rect 345020 132336 345072 132388
rect 252376 131520 252428 131572
rect 260288 131520 260340 131572
rect 294788 131248 294840 131300
rect 307668 131248 307720 131300
rect 207664 131180 207716 131232
rect 213920 131180 213972 131232
rect 278044 131180 278096 131232
rect 307392 131180 307444 131232
rect 189724 131112 189776 131164
rect 214012 131112 214064 131164
rect 271144 131112 271196 131164
rect 307576 131112 307628 131164
rect 252284 131044 252336 131096
rect 291844 131044 291896 131096
rect 324412 131044 324464 131096
rect 342444 131044 342496 131096
rect 252468 130976 252520 131028
rect 267280 130976 267332 131028
rect 324320 130976 324372 131028
rect 331220 130976 331272 131028
rect 252376 130364 252428 130416
rect 261576 130364 261628 130416
rect 296260 129888 296312 129940
rect 307668 129888 307720 129940
rect 199384 129820 199436 129872
rect 214012 129820 214064 129872
rect 285128 129820 285180 129872
rect 307484 129820 307536 129872
rect 171876 129752 171928 129804
rect 213920 129752 213972 129804
rect 273996 129752 274048 129804
rect 307576 129752 307628 129804
rect 252468 129684 252520 129736
rect 269856 129684 269908 129736
rect 324412 129684 324464 129736
rect 346584 129684 346636 129736
rect 252284 129616 252336 129668
rect 261668 129616 261720 129668
rect 324320 129616 324372 129668
rect 330116 129616 330168 129668
rect 252008 129004 252060 129056
rect 305736 129004 305788 129056
rect 301596 128460 301648 128512
rect 306748 128460 306800 128512
rect 296076 128392 296128 128444
rect 307668 128392 307720 128444
rect 178776 128324 178828 128376
rect 213920 128324 213972 128376
rect 276664 128324 276716 128376
rect 307576 128324 307628 128376
rect 252376 128256 252428 128308
rect 282276 128256 282328 128308
rect 324320 128256 324372 128308
rect 328552 128256 328604 128308
rect 252468 128188 252520 128240
rect 271328 128188 271380 128240
rect 252468 127440 252520 127492
rect 258908 127440 258960 127492
rect 289176 127100 289228 127152
rect 307668 127100 307720 127152
rect 272524 127032 272576 127084
rect 307576 127032 307628 127084
rect 271236 126964 271288 127016
rect 307484 126964 307536 127016
rect 252468 126896 252520 126948
rect 272616 126896 272668 126948
rect 324320 126896 324372 126948
rect 328460 126896 328512 126948
rect 392584 126896 392636 126948
rect 580172 126896 580224 126948
rect 252376 126624 252428 126676
rect 258816 126624 258868 126676
rect 252192 126216 252244 126268
rect 300400 126216 300452 126268
rect 300124 125740 300176 125792
rect 307668 125740 307720 125792
rect 191196 125672 191248 125724
rect 214012 125672 214064 125724
rect 286508 125672 286560 125724
rect 307576 125672 307628 125724
rect 62028 125604 62080 125656
rect 65156 125604 65208 125656
rect 169116 125604 169168 125656
rect 213920 125604 213972 125656
rect 273904 125604 273956 125656
rect 307484 125604 307536 125656
rect 252468 125536 252520 125588
rect 274088 125536 274140 125588
rect 252376 125468 252428 125520
rect 253480 125468 253532 125520
rect 275376 124924 275428 124976
rect 307300 124924 307352 124976
rect 252284 124856 252336 124908
rect 297456 124856 297508 124908
rect 303068 124312 303120 124364
rect 306932 124312 306984 124364
rect 180064 124244 180116 124296
rect 213920 124244 213972 124296
rect 298928 124244 298980 124296
rect 307576 124244 307628 124296
rect 170588 124176 170640 124228
rect 214012 124176 214064 124228
rect 295984 124176 296036 124228
rect 307668 124176 307720 124228
rect 252468 124108 252520 124160
rect 269764 124108 269816 124160
rect 324320 124108 324372 124160
rect 340880 124108 340932 124160
rect 252376 124040 252428 124092
rect 261484 124040 261536 124092
rect 252284 123428 252336 123480
rect 304540 123428 304592 123480
rect 211804 123360 211856 123412
rect 213920 123360 213972 123412
rect 304356 122952 304408 123004
rect 307668 122952 307720 123004
rect 292028 122884 292080 122936
rect 307484 122884 307536 122936
rect 195336 122816 195388 122868
rect 213920 122816 213972 122868
rect 282368 122816 282420 122868
rect 307576 122816 307628 122868
rect 324320 122748 324372 122800
rect 336740 122748 336792 122800
rect 252376 122680 252428 122732
rect 286324 122680 286376 122732
rect 252468 122612 252520 122664
rect 289360 122612 289412 122664
rect 297548 121592 297600 121644
rect 307576 121592 307628 121644
rect 202236 121524 202288 121576
rect 213920 121524 213972 121576
rect 289268 121524 289320 121576
rect 307668 121524 307720 121576
rect 182824 121456 182876 121508
rect 214012 121456 214064 121508
rect 286416 121456 286468 121508
rect 307484 121456 307536 121508
rect 252376 121388 252428 121440
rect 290648 121388 290700 121440
rect 324412 121388 324464 121440
rect 343824 121388 343876 121440
rect 324320 121320 324372 121372
rect 338304 121320 338356 121372
rect 251916 120708 251968 120760
rect 268476 120708 268528 120760
rect 252468 120640 252520 120692
rect 260104 120640 260156 120692
rect 291844 120232 291896 120284
rect 307668 120232 307720 120284
rect 290464 120164 290516 120216
rect 307576 120164 307628 120216
rect 170680 120096 170732 120148
rect 213920 120096 213972 120148
rect 269764 120096 269816 120148
rect 307484 120096 307536 120148
rect 252376 120028 252428 120080
rect 298744 120028 298796 120080
rect 324320 120028 324372 120080
rect 338212 120028 338264 120080
rect 252468 119960 252520 120012
rect 262956 119960 263008 120012
rect 252468 119416 252520 119468
rect 258724 119416 258776 119468
rect 263048 119348 263100 119400
rect 307392 119348 307444 119400
rect 178868 118804 178920 118856
rect 214012 118804 214064 118856
rect 298836 118804 298888 118856
rect 307668 118804 307720 118856
rect 172060 118736 172112 118788
rect 214104 118736 214156 118788
rect 167920 118668 167972 118720
rect 213920 118668 213972 118720
rect 301688 118668 301740 118720
rect 307484 118668 307536 118720
rect 252468 118600 252520 118652
rect 267096 118600 267148 118652
rect 324320 118600 324372 118652
rect 340972 118600 341024 118652
rect 252376 118532 252428 118584
rect 256148 118532 256200 118584
rect 324412 118532 324464 118584
rect 332692 118532 332744 118584
rect 174728 117920 174780 117972
rect 214748 117920 214800 117972
rect 252284 117920 252336 117972
rect 296168 117920 296220 117972
rect 293316 117444 293368 117496
rect 307668 117444 307720 117496
rect 268384 117376 268436 117428
rect 307576 117376 307628 117428
rect 181444 117308 181496 117360
rect 213920 117308 213972 117360
rect 260104 117308 260156 117360
rect 306564 117308 306616 117360
rect 252468 117240 252520 117292
rect 262864 117240 262916 117292
rect 324320 117240 324372 117292
rect 333980 117240 334032 117292
rect 252100 116560 252152 116612
rect 281080 116560 281132 116612
rect 252468 116084 252520 116136
rect 260196 116084 260248 116136
rect 296168 116084 296220 116136
rect 307576 116084 307628 116136
rect 186964 116016 187016 116068
rect 213920 116016 213972 116068
rect 280896 116016 280948 116068
rect 307668 116016 307720 116068
rect 176108 115948 176160 116000
rect 214012 115948 214064 116000
rect 267188 115948 267240 116000
rect 306748 115948 306800 116000
rect 252376 115880 252428 115932
rect 264520 115880 264572 115932
rect 252284 115200 252336 115252
rect 282460 115200 282512 115252
rect 293408 114656 293460 114708
rect 307576 114656 307628 114708
rect 180156 114588 180208 114640
rect 213920 114588 213972 114640
rect 287888 114588 287940 114640
rect 307668 114588 307720 114640
rect 176016 114520 176068 114572
rect 214012 114520 214064 114572
rect 264244 114520 264296 114572
rect 307484 114520 307536 114572
rect 252468 114452 252520 114504
rect 300216 114452 300268 114504
rect 324320 114452 324372 114504
rect 342352 114452 342404 114504
rect 252376 114384 252428 114436
rect 285036 114384 285088 114436
rect 324412 114384 324464 114436
rect 335544 114384 335596 114436
rect 211896 113228 211948 113280
rect 214012 113228 214064 113280
rect 294604 113228 294656 113280
rect 307668 113228 307720 113280
rect 198096 113160 198148 113212
rect 213920 113160 213972 113212
rect 284944 113160 284996 113212
rect 307576 113160 307628 113212
rect 252468 113092 252520 113144
rect 299112 113092 299164 113144
rect 324320 113092 324372 113144
rect 337016 113092 337068 113144
rect 252008 112412 252060 112464
rect 305644 112412 305696 112464
rect 204996 111868 205048 111920
rect 214012 111868 214064 111920
rect 301504 111868 301556 111920
rect 307484 111868 307536 111920
rect 169208 111800 169260 111852
rect 213920 111800 213972 111852
rect 253204 111800 253256 111852
rect 307668 111800 307720 111852
rect 3148 111732 3200 111784
rect 17224 111732 17276 111784
rect 168012 111732 168064 111784
rect 171968 111732 172020 111784
rect 252468 111732 252520 111784
rect 304264 111732 304316 111784
rect 252376 111664 252428 111716
rect 256056 111664 256108 111716
rect 252284 111052 252336 111104
rect 301780 111052 301832 111104
rect 192484 110508 192536 110560
rect 214012 110508 214064 110560
rect 300216 110508 300268 110560
rect 307576 110508 307628 110560
rect 173440 110440 173492 110492
rect 213920 110440 213972 110492
rect 303160 110440 303212 110492
rect 307668 110440 307720 110492
rect 168104 110372 168156 110424
rect 175924 110372 175976 110424
rect 252376 110372 252428 110424
rect 287980 110372 288032 110424
rect 252468 110304 252520 110356
rect 264336 110304 264388 110356
rect 251640 110236 251692 110288
rect 254584 110236 254636 110288
rect 304540 109148 304592 109200
rect 307484 109148 307536 109200
rect 209136 109080 209188 109132
rect 214012 109080 214064 109132
rect 287796 109080 287848 109132
rect 307576 109080 307628 109132
rect 174636 109012 174688 109064
rect 213920 109012 213972 109064
rect 262864 109012 262916 109064
rect 307668 109012 307720 109064
rect 168012 108944 168064 108996
rect 177580 108944 177632 108996
rect 252376 108944 252428 108996
rect 292120 108944 292172 108996
rect 324320 108944 324372 108996
rect 353300 108944 353352 108996
rect 252468 108876 252520 108928
rect 275376 108876 275428 108928
rect 282276 107856 282328 107908
rect 307668 107856 307720 107908
rect 292212 107720 292264 107772
rect 307668 107720 307720 107772
rect 177672 107652 177724 107704
rect 213920 107652 213972 107704
rect 302976 107652 303028 107704
rect 307576 107652 307628 107704
rect 252376 107584 252428 107636
rect 305920 107584 305972 107636
rect 252468 107516 252520 107568
rect 264428 107516 264480 107568
rect 252192 107448 252244 107500
rect 254676 107448 254728 107500
rect 268476 106428 268528 106480
rect 307484 106428 307536 106480
rect 304264 106360 304316 106412
rect 307668 106360 307720 106412
rect 169300 106292 169352 106344
rect 213920 106292 213972 106344
rect 252468 106224 252520 106276
rect 285220 106224 285272 106276
rect 252284 106156 252336 106208
rect 255964 106156 256016 106208
rect 252376 105544 252428 105596
rect 299020 105544 299072 105596
rect 300492 105000 300544 105052
rect 307668 105000 307720 105052
rect 207756 104932 207808 104984
rect 213920 104932 213972 104984
rect 298744 104932 298796 104984
rect 307484 104932 307536 104984
rect 199476 104864 199528 104916
rect 214012 104864 214064 104916
rect 285036 104864 285088 104916
rect 307576 104864 307628 104916
rect 252468 104796 252520 104848
rect 265624 104796 265676 104848
rect 252284 104728 252336 104780
rect 257436 104728 257488 104780
rect 251272 104116 251324 104168
rect 275284 104116 275336 104168
rect 210608 103844 210660 103896
rect 213920 103844 213972 103896
rect 279424 103572 279476 103624
rect 307668 103572 307720 103624
rect 171968 103504 172020 103556
rect 213920 103504 213972 103556
rect 267096 103504 267148 103556
rect 307576 103504 307628 103556
rect 252468 103436 252520 103488
rect 268568 103436 268620 103488
rect 324412 103436 324464 103488
rect 339684 103436 339736 103488
rect 251180 103300 251232 103352
rect 253388 103300 253440 103352
rect 252192 102756 252244 102808
rect 269948 102756 270000 102808
rect 294696 102280 294748 102332
rect 306932 102280 306984 102332
rect 275284 102212 275336 102264
rect 307576 102212 307628 102264
rect 269856 102144 269908 102196
rect 307668 102144 307720 102196
rect 251364 102076 251416 102128
rect 253296 102076 253348 102128
rect 252468 102008 252520 102060
rect 280988 102008 281040 102060
rect 252284 101396 252336 101448
rect 300308 101396 300360 101448
rect 300400 100852 300452 100904
rect 307576 100852 307628 100904
rect 299020 100784 299072 100836
rect 307484 100784 307536 100836
rect 283656 100716 283708 100768
rect 307668 100716 307720 100768
rect 252376 100648 252428 100700
rect 304448 100648 304500 100700
rect 252468 100580 252520 100632
rect 294880 100580 294932 100632
rect 166540 99424 166592 99476
rect 213920 99424 213972 99476
rect 297456 99424 297508 99476
rect 307576 99424 307628 99476
rect 166356 99356 166408 99408
rect 214012 99356 214064 99408
rect 290648 99356 290700 99408
rect 307668 99356 307720 99408
rect 252376 99288 252428 99340
rect 286600 99288 286652 99340
rect 252468 99220 252520 99272
rect 257344 99220 257396 99272
rect 166448 98064 166500 98116
rect 214012 98064 214064 98116
rect 286324 98064 286376 98116
rect 307576 98064 307628 98116
rect 164976 97996 165028 98048
rect 213920 97996 213972 98048
rect 258724 97996 258776 98048
rect 307668 97996 307720 98048
rect 252468 97928 252520 97980
rect 263048 97928 263100 97980
rect 2780 97724 2832 97776
rect 4804 97724 4856 97776
rect 289360 96704 289412 96756
rect 306932 96704 306984 96756
rect 210516 96636 210568 96688
rect 213920 96636 213972 96688
rect 255964 96636 256016 96688
rect 307668 96636 307720 96688
rect 308496 96568 308548 96620
rect 321468 96568 321520 96620
rect 198188 95208 198240 95260
rect 213920 95208 213972 95260
rect 249064 95208 249116 95260
rect 307668 95208 307720 95260
rect 196624 95140 196676 95192
rect 324320 95140 324372 95192
rect 308404 95072 308456 95124
rect 324412 95072 324464 95124
rect 309784 95004 309836 95056
rect 321376 95004 321428 95056
rect 122840 94460 122892 94512
rect 214840 94460 214892 94512
rect 151636 94052 151688 94104
rect 178684 94052 178736 94104
rect 129372 93984 129424 94036
rect 166264 93984 166316 94036
rect 111984 93916 112036 93968
rect 170496 93916 170548 93968
rect 113732 93848 113784 93900
rect 172060 93848 172112 93900
rect 62028 93780 62080 93832
rect 210608 93780 210660 93832
rect 216036 93780 216088 93832
rect 321652 93780 321704 93832
rect 188344 93712 188396 93764
rect 324504 93712 324556 93764
rect 191104 93644 191156 93696
rect 321560 93644 321612 93696
rect 133144 93372 133196 93424
rect 174544 93372 174596 93424
rect 118056 93304 118108 93356
rect 170404 93304 170456 93356
rect 120632 93236 120684 93288
rect 195336 93236 195388 93288
rect 107752 93168 107804 93220
rect 186964 93168 187016 93220
rect 85672 93100 85724 93152
rect 164976 93100 165028 93152
rect 115480 92420 115532 92472
rect 204904 92420 204956 92472
rect 95056 92352 95108 92404
rect 122840 92352 122892 92404
rect 125968 92352 126020 92404
rect 206376 92352 206428 92404
rect 116768 92284 116820 92336
rect 174728 92284 174780 92336
rect 151728 92216 151780 92268
rect 198004 92216 198056 92268
rect 130752 92148 130804 92200
rect 169024 92148 169076 92200
rect 152096 92080 152148 92132
rect 173256 92080 173308 92132
rect 238024 91808 238076 91860
rect 251180 91808 251232 91860
rect 206284 91740 206336 91792
rect 307300 91740 307352 91792
rect 91652 91128 91704 91180
rect 108304 91128 108356 91180
rect 85120 91060 85172 91112
rect 129004 91060 129056 91112
rect 66076 90992 66128 91044
rect 171968 90992 172020 91044
rect 120540 90924 120592 90976
rect 209044 90924 209096 90976
rect 106004 90856 106056 90908
rect 189724 90856 189776 90908
rect 110328 90788 110380 90840
rect 176108 90788 176160 90840
rect 125508 90720 125560 90772
rect 169116 90720 169168 90772
rect 136456 90652 136508 90704
rect 167736 90652 167788 90704
rect 177304 90312 177356 90364
rect 307208 90312 307260 90364
rect 64788 89632 64840 89684
rect 216220 89632 216272 89684
rect 90640 89564 90692 89616
rect 199476 89564 199528 89616
rect 102692 89496 102744 89548
rect 211896 89496 211948 89548
rect 100024 89428 100076 89480
rect 192484 89428 192536 89480
rect 115388 89360 115440 89412
rect 178868 89360 178920 89412
rect 151268 89292 151320 89344
rect 213184 89292 213236 89344
rect 215944 88952 215996 89004
rect 307116 88952 307168 89004
rect 67640 88272 67692 88324
rect 214932 88272 214984 88324
rect 67456 88204 67508 88256
rect 214564 88204 214616 88256
rect 126520 88136 126572 88188
rect 191196 88136 191248 88188
rect 111248 88068 111300 88120
rect 167828 88068 167880 88120
rect 117136 88000 117188 88052
rect 170680 88000 170732 88052
rect 123484 87932 123536 87984
rect 177396 87932 177448 87984
rect 101864 86912 101916 86964
rect 204996 86912 205048 86964
rect 88064 86844 88116 86896
rect 166540 86844 166592 86896
rect 134616 86776 134668 86828
rect 210424 86776 210476 86828
rect 109592 86708 109644 86760
rect 177488 86708 177540 86760
rect 112352 86640 112404 86692
rect 167920 86640 167972 86692
rect 124128 86572 124180 86624
rect 170588 86572 170640 86624
rect 3516 85484 3568 85536
rect 22744 85484 22796 85536
rect 67364 85484 67416 85536
rect 210516 85484 210568 85536
rect 111432 85416 111484 85468
rect 213368 85416 213420 85468
rect 104256 85348 104308 85400
rect 198096 85348 198148 85400
rect 100576 85280 100628 85332
rect 169208 85280 169260 85332
rect 122840 85212 122892 85264
rect 180064 85212 180116 85264
rect 132408 85144 132460 85196
rect 173164 85144 173216 85196
rect 104808 84124 104860 84176
rect 207664 84124 207716 84176
rect 118608 84056 118660 84108
rect 202236 84056 202288 84108
rect 86868 83988 86920 84040
rect 166448 83988 166500 84040
rect 96528 83920 96580 83972
rect 174636 83920 174688 83972
rect 106188 83852 106240 83904
rect 180156 83852 180208 83904
rect 122656 83784 122708 83836
rect 171784 83784 171836 83836
rect 122748 82764 122800 82816
rect 211804 82764 211856 82816
rect 89628 82696 89680 82748
rect 166356 82696 166408 82748
rect 99104 82628 99156 82680
rect 173440 82628 173492 82680
rect 110144 82560 110196 82612
rect 181444 82560 181496 82612
rect 101956 82492 102008 82544
rect 171876 82492 171928 82544
rect 125416 82424 125468 82476
rect 167644 82424 167696 82476
rect 108304 81336 108356 81388
rect 214656 81336 214708 81388
rect 93768 81268 93820 81320
rect 169300 81268 169352 81320
rect 128268 81200 128320 81252
rect 202144 81200 202196 81252
rect 107476 81132 107528 81184
rect 173348 81132 173400 81184
rect 115848 79976 115900 80028
rect 213276 79976 213328 80028
rect 108948 79908 109000 79960
rect 196716 79908 196768 79960
rect 95148 79840 95200 79892
rect 177672 79840 177724 79892
rect 114468 79772 114520 79824
rect 195244 79772 195296 79824
rect 97908 78616 97960 78668
rect 209136 78616 209188 78668
rect 129004 78548 129056 78600
rect 216128 78548 216180 78600
rect 102048 78480 102100 78532
rect 178776 78480 178828 78532
rect 119988 78412 120040 78464
rect 182824 78412 182876 78464
rect 75828 77188 75880 77240
rect 198188 77188 198240 77240
rect 124220 76576 124272 76628
rect 279516 76576 279568 76628
rect 82820 76508 82872 76560
rect 292212 76508 292264 76560
rect 107568 75828 107620 75880
rect 176016 75828 176068 75880
rect 115940 75216 115992 75268
rect 303068 75216 303120 75268
rect 23480 75148 23532 75200
rect 272524 75148 272576 75200
rect 93860 73856 93912 73908
rect 306012 73856 306064 73908
rect 56600 73788 56652 73840
rect 294788 73788 294840 73840
rect 118700 72496 118752 72548
rect 298928 72496 298980 72548
rect 64880 72428 64932 72480
rect 300492 72428 300544 72480
rect 3516 71680 3568 71732
rect 53104 71680 53156 71732
rect 103520 71068 103572 71120
rect 304540 71068 304592 71120
rect 52460 71000 52512 71052
rect 296260 71000 296312 71052
rect 9680 69640 9732 69692
rect 286508 69640 286560 69692
rect 110420 68348 110472 68400
rect 303160 68348 303212 68400
rect 44180 68280 44232 68332
rect 267188 68280 267240 68332
rect 114560 66920 114612 66972
rect 300216 66920 300268 66972
rect 34520 66852 34572 66904
rect 293408 66852 293460 66904
rect 121460 65560 121512 65612
rect 253204 65560 253256 65612
rect 30380 65492 30432 65544
rect 287888 65492 287940 65544
rect 69020 64200 69072 64252
rect 305828 64200 305880 64252
rect 29000 64132 29052 64184
rect 300400 64132 300452 64184
rect 71780 62772 71832 62824
rect 268476 62772 268528 62824
rect 98000 61344 98052 61396
rect 282368 61344 282420 61396
rect 184204 60664 184256 60716
rect 580172 60664 580224 60716
rect 4160 59984 4212 60036
rect 249064 59984 249116 60036
rect 70400 58692 70452 58744
rect 290556 58692 290608 58744
rect 33140 58624 33192 58676
rect 299020 58624 299072 58676
rect 85580 57196 85632 57248
rect 291936 57196 291988 57248
rect 45560 55904 45612 55956
rect 273996 55904 274048 55956
rect 73160 55836 73212 55888
rect 301688 55836 301740 55888
rect 86960 53116 87012 53168
rect 289268 53116 289320 53168
rect 27620 53048 27672 53100
rect 271236 53048 271288 53100
rect 91100 51756 91152 51808
rect 297548 51756 297600 51808
rect 19340 51688 19392 51740
rect 289176 51688 289228 51740
rect 104900 50396 104952 50448
rect 292028 50396 292080 50448
rect 81440 50328 81492 50380
rect 276756 50328 276808 50380
rect 102140 49036 102192 49088
rect 304356 49036 304408 49088
rect 60740 48968 60792 49020
rect 271144 48968 271196 49020
rect 88340 47540 88392 47592
rect 278136 47540 278188 47592
rect 20 46860 72 46912
rect 1308 46860 1360 46912
rect 249156 46860 249208 46912
rect 122840 46180 122892 46232
rect 300124 46180 300176 46232
rect 3424 45500 3476 45552
rect 15844 45500 15896 45552
rect 93952 44888 94004 44940
rect 286416 44888 286468 44940
rect 13820 44820 13872 44872
rect 273904 44820 273956 44872
rect 84200 43460 84252 43512
rect 269764 43460 269816 43512
rect 95240 43392 95292 43444
rect 287704 43392 287756 43444
rect 80060 42100 80112 42152
rect 290464 42100 290516 42152
rect 35992 42032 36044 42084
rect 301596 42032 301648 42084
rect 77300 40740 77352 40792
rect 291844 40740 291896 40792
rect 42800 40672 42852 40724
rect 285128 40672 285180 40724
rect 57980 39380 58032 39432
rect 267096 39380 267148 39432
rect 66260 39312 66312 39364
rect 298836 39312 298888 39364
rect 99380 37952 99432 38004
rect 283564 37952 283616 38004
rect 24860 37884 24912 37936
rect 307024 37884 307076 37936
rect 92480 36592 92532 36644
rect 302884 36592 302936 36644
rect 16580 36524 16632 36576
rect 290648 36524 290700 36576
rect 40040 35232 40092 35284
rect 269856 35232 269908 35284
rect 52552 35164 52604 35216
rect 293316 35164 293368 35216
rect 106280 33804 106332 33856
rect 293224 33804 293276 33856
rect 48320 33736 48372 33788
rect 296168 33736 296220 33788
rect 3148 33056 3200 33108
rect 32404 33056 32456 33108
rect 2780 31016 2832 31068
rect 289360 31016 289412 31068
rect 44272 29588 44324 29640
rect 294696 29588 294748 29640
rect 75920 28296 75972 28348
rect 305736 28296 305788 28348
rect 26240 28228 26292 28280
rect 283656 28228 283708 28280
rect 96620 26936 96672 26988
rect 262864 26936 262916 26988
rect 20720 26868 20772 26920
rect 297456 26868 297508 26920
rect 118792 25576 118844 25628
rect 301504 25576 301556 25628
rect 37280 25508 37332 25560
rect 264244 25508 264296 25560
rect 107660 24148 107712 24200
rect 305644 24148 305696 24200
rect 41420 24080 41472 24132
rect 280896 24080 280948 24132
rect 100760 22788 100812 22840
rect 287796 22788 287848 22840
rect 63500 22720 63552 22772
rect 278044 22720 278096 22772
rect 85672 21428 85724 21480
rect 302976 21428 303028 21480
rect 31760 21360 31812 21412
rect 296076 21360 296128 21412
rect 3424 20612 3476 20664
rect 11704 20612 11756 20664
rect 17960 19932 18012 19984
rect 294604 19932 294656 19984
rect 89720 18572 89772 18624
rect 282276 18572 282328 18624
rect 78680 17280 78732 17332
rect 304264 17280 304316 17332
rect 38660 17212 38712 17264
rect 276664 17212 276716 17264
rect 69112 15920 69164 15972
rect 298744 15920 298796 15972
rect 11152 15852 11204 15904
rect 255964 15852 256016 15904
rect 61568 14492 61620 14544
rect 285036 14492 285088 14544
rect 20168 14424 20220 14476
rect 258724 14424 258776 14476
rect 3424 13132 3476 13184
rect 51724 13132 51776 13184
rect 51080 13064 51132 13116
rect 279424 13064 279476 13116
rect 120632 11772 120684 11824
rect 250444 11772 250496 11824
rect 7656 11704 7708 11756
rect 286324 11704 286376 11756
rect 117320 10344 117372 10396
rect 267004 10344 267056 10396
rect 2872 10276 2924 10328
rect 289084 10276 289136 10328
rect 7472 9596 7524 9648
rect 8208 9596 8260 9648
rect 251180 9596 251232 9648
rect 75000 8916 75052 8968
rect 282184 8916 282236 8968
rect 1676 8304 1728 8356
rect 7472 8304 7524 8356
rect 103336 7624 103388 7676
rect 297364 7624 297416 7676
rect 47860 7556 47912 7608
rect 275284 7556 275336 7608
rect 27712 6128 27764 6180
rect 284944 6128 284996 6180
rect 56048 4768 56100 4820
rect 268384 4768 268436 4820
rect 125876 3680 125928 3732
rect 164884 3680 164936 3732
rect 110512 3612 110564 3664
rect 67916 3544 67968 3596
rect 2780 3476 2832 3528
rect 3700 3476 3752 3528
rect 11060 3476 11112 3528
rect 11980 3476 12032 3528
rect 35900 3476 35952 3528
rect 36820 3476 36872 3528
rect 44180 3476 44232 3528
rect 45100 3476 45152 3528
rect 52460 3476 52512 3528
rect 53380 3476 53432 3528
rect 69020 3476 69072 3528
rect 69940 3476 69992 3528
rect 110420 3544 110472 3596
rect 111616 3544 111668 3596
rect 112812 3612 112864 3664
rect 206284 3612 206336 3664
rect 215944 3544 215996 3596
rect 177304 3476 177356 3528
rect 235816 3476 235868 3528
rect 238024 3476 238076 3528
rect 23020 3408 23072 3460
rect 47584 3408 47636 3460
rect 63224 3408 63276 3460
rect 260104 3408 260156 3460
rect 118700 3340 118752 3392
rect 119896 3340 119948 3392
rect 114008 2116 114060 2168
rect 280804 2116 280856 2168
rect 109316 2048 109368 2100
rect 295984 2048 296036 2100
<< metal2 >>
rect 6932 703582 7972 703610
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3238 566944 3294 566953
rect 3238 566879 3294 566888
rect 3252 565894 3280 566879
rect 3240 565888 3292 565894
rect 3240 565830 3292 565836
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2976 527202 3004 527847
rect 2964 527196 3016 527202
rect 2964 527138 3016 527144
rect 3330 501800 3386 501809
rect 3330 501735 3386 501744
rect 3344 501022 3372 501735
rect 3332 501016 3384 501022
rect 3332 500958 3384 500964
rect 3054 475688 3110 475697
rect 3054 475623 3110 475632
rect 3068 474774 3096 475623
rect 3056 474768 3108 474774
rect 3056 474710 3108 474716
rect 3330 462632 3386 462641
rect 3330 462567 3386 462576
rect 3344 462398 3372 462567
rect 3332 462392 3384 462398
rect 3332 462334 3384 462340
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 3344 448594 3372 449511
rect 3332 448588 3384 448594
rect 3332 448530 3384 448536
rect 2778 423600 2834 423609
rect 2778 423535 2780 423544
rect 2832 423535 2834 423544
rect 2780 423506 2832 423512
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3344 409902 3372 410479
rect 3332 409896 3384 409902
rect 3332 409838 3384 409844
rect 3332 397520 3384 397526
rect 3330 397488 3332 397497
rect 3384 397488 3386 397497
rect 3330 397423 3386 397432
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3344 371278 3372 371311
rect 3332 371272 3384 371278
rect 3332 371214 3384 371220
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3344 357474 3372 358391
rect 3332 357468 3384 357474
rect 3332 357410 3384 357416
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3436 324970 3464 684247
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3528 656946 3556 658135
rect 3516 656940 3568 656946
rect 3516 656882 3568 656888
rect 3516 632120 3568 632126
rect 3514 632088 3516 632097
rect 3568 632088 3570 632097
rect 3514 632023 3570 632032
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618322 3556 619103
rect 3516 618316 3568 618322
rect 3516 618258 3568 618264
rect 3514 606112 3570 606121
rect 3514 606047 3570 606056
rect 3528 605878 3556 606047
rect 3516 605872 3568 605878
rect 3516 605814 3568 605820
rect 3514 514856 3570 514865
rect 3514 514791 3570 514800
rect 3424 324964 3476 324970
rect 3424 324906 3476 324912
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3344 318850 3372 319223
rect 3332 318844 3384 318850
rect 3332 318786 3384 318792
rect 3528 315314 3556 514791
rect 4804 423564 4856 423570
rect 4804 423506 4856 423512
rect 3516 315308 3568 315314
rect 3516 315250 3568 315256
rect 3238 306232 3294 306241
rect 3238 306167 3294 306176
rect 3252 305046 3280 306167
rect 3240 305040 3292 305046
rect 3240 304982 3292 304988
rect 4816 298790 4844 423506
rect 4804 298784 4856 298790
rect 4804 298726 4856 298732
rect 3424 294092 3476 294098
rect 3424 294034 3476 294040
rect 2778 293176 2834 293185
rect 2778 293111 2834 293120
rect 2792 292874 2820 293111
rect 2780 292868 2832 292874
rect 2780 292810 2832 292816
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3160 253978 3188 254079
rect 3148 253972 3200 253978
rect 3148 253914 3200 253920
rect 3054 241088 3110 241097
rect 3054 241023 3110 241032
rect 3068 240174 3096 241023
rect 3056 240168 3108 240174
rect 3056 240110 3108 240116
rect 1308 220244 1360 220250
rect 1308 220186 1360 220192
rect 1320 46918 1348 220186
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3056 202836 3108 202842
rect 3056 202778 3108 202784
rect 3068 201929 3096 202778
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 2780 97776 2832 97782
rect 2780 97718 2832 97724
rect 2792 97617 2820 97718
rect 2778 97608 2834 97617
rect 2778 97543 2834 97552
rect 3436 58585 3464 294034
rect 4804 292868 4856 292874
rect 4804 292810 4856 292816
rect 3516 291848 3568 291854
rect 3516 291790 3568 291796
rect 3528 188873 3556 291790
rect 3606 267200 3662 267209
rect 3606 267135 3662 267144
rect 3620 239426 3648 267135
rect 4816 244254 4844 292810
rect 6932 269822 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 24320 699718 24348 703520
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 25504 699712 25556 699718
rect 25504 699654 25556 699660
rect 15844 656940 15896 656946
rect 15844 656882 15896 656888
rect 14464 605872 14516 605878
rect 14464 605814 14516 605820
rect 11704 318844 11756 318850
rect 11704 318786 11756 318792
rect 11716 318102 11744 318786
rect 11704 318096 11756 318102
rect 11704 318038 11756 318044
rect 14476 311166 14504 605814
rect 14464 311160 14516 311166
rect 14464 311102 14516 311108
rect 15856 309806 15884 656882
rect 21364 632120 21416 632126
rect 21364 632062 21416 632068
rect 17224 618316 17276 618322
rect 17224 618258 17276 618264
rect 15844 309800 15896 309806
rect 15844 309742 15896 309748
rect 11704 295656 11756 295662
rect 11704 295598 11756 295604
rect 8208 292868 8260 292874
rect 8208 292810 8260 292816
rect 6920 269816 6972 269822
rect 6920 269758 6972 269764
rect 4804 244248 4856 244254
rect 4804 244190 4856 244196
rect 3608 239420 3660 239426
rect 3608 239362 3660 239368
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 4804 177336 4856 177342
rect 4804 177278 4856 177284
rect 3516 150408 3568 150414
rect 3516 150350 3568 150356
rect 3528 149841 3556 150350
rect 3514 149832 3570 149841
rect 3514 149767 3570 149776
rect 3516 137964 3568 137970
rect 3516 137906 3568 137912
rect 3528 136785 3556 137906
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 4816 97782 4844 177278
rect 4804 97776 4856 97782
rect 4804 97718 4856 97724
rect 3516 85536 3568 85542
rect 3516 85478 3568 85484
rect 3528 84697 3556 85478
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 3516 71732 3568 71738
rect 3516 71674 3568 71680
rect 3528 71641 3556 71674
rect 3514 71632 3570 71641
rect 3514 71567 3570 71576
rect 4160 60036 4212 60042
rect 4160 59978 4212 59984
rect 3422 58576 3478 58585
rect 3422 58511 3478 58520
rect 20 46912 72 46918
rect 20 46854 72 46860
rect 1308 46912 1360 46918
rect 1308 46854 1360 46860
rect 32 16574 60 46854
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3148 33108 3200 33114
rect 3148 33050 3200 33056
rect 3160 32473 3188 33050
rect 3146 32464 3202 32473
rect 3146 32399 3202 32408
rect 2780 31068 2832 31074
rect 2780 31010 2832 31016
rect 32 16546 152 16574
rect 124 354 152 16546
rect 1676 8356 1728 8362
rect 1676 8298 1728 8304
rect 1688 480 1716 8298
rect 2792 3534 2820 31010
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4172 16574 4200 59978
rect 4172 16546 5304 16574
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 2872 10328 2924 10334
rect 2872 10270 2924 10276
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2884 480 2912 10270
rect 3436 6497 3464 13126
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 542 354 654 480
rect 124 326 654 354
rect 542 -960 654 326
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3712 354 3740 3470
rect 5276 480 5304 16546
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 7472 9648 7524 9654
rect 7472 9590 7524 9596
rect 7484 8362 7512 9590
rect 7472 8356 7524 8362
rect 7472 8298 7524 8304
rect 6458 4856 6514 4865
rect 6458 4791 6514 4800
rect 6472 480 6500 4791
rect 7668 480 7696 11698
rect 8220 9654 8248 292810
rect 9680 69692 9732 69698
rect 9680 69634 9732 69640
rect 8298 61432 8354 61441
rect 8298 61367 8354 61376
rect 8312 16574 8340 61367
rect 8312 16546 8800 16574
rect 8208 9648 8260 9654
rect 8208 9590 8260 9596
rect 8772 480 8800 16546
rect 4038 354 4150 480
rect 3712 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 69634
rect 11716 20670 11744 295598
rect 17236 274650 17264 618258
rect 18604 553444 18656 553450
rect 18604 553386 18656 553392
rect 17224 274644 17276 274650
rect 17224 274586 17276 274592
rect 17224 263628 17276 263634
rect 17224 263570 17276 263576
rect 14464 256760 14516 256766
rect 14464 256702 14516 256708
rect 14476 137970 14504 256702
rect 15200 240168 15252 240174
rect 15200 240110 15252 240116
rect 15212 238746 15240 240110
rect 15200 238740 15252 238746
rect 15200 238682 15252 238688
rect 15844 231192 15896 231198
rect 15844 231134 15896 231140
rect 14464 137964 14516 137970
rect 14464 137906 14516 137912
rect 15198 57216 15254 57225
rect 15198 57151 15254 57160
rect 12438 54496 12494 54505
rect 12438 54431 12494 54440
rect 11704 20664 11756 20670
rect 11704 20606 11756 20612
rect 11058 18592 11114 18601
rect 11058 18527 11114 18536
rect 11072 3534 11100 18527
rect 12452 16574 12480 54431
rect 13820 44872 13872 44878
rect 13820 44814 13872 44820
rect 13832 16574 13860 44814
rect 15212 16574 15240 57151
rect 15856 45558 15884 231134
rect 17236 215286 17264 263570
rect 18616 263566 18644 553386
rect 21376 266354 21404 632062
rect 22744 448588 22796 448594
rect 22744 448530 22796 448536
rect 22756 301510 22784 448530
rect 25516 304298 25544 699654
rect 32404 670744 32456 670750
rect 32404 670686 32456 670692
rect 29644 565888 29696 565894
rect 29644 565830 29696 565836
rect 25504 304292 25556 304298
rect 25504 304234 25556 304240
rect 22744 301504 22796 301510
rect 22744 301446 22796 301452
rect 25504 289876 25556 289882
rect 25504 289818 25556 289824
rect 21364 266348 21416 266354
rect 21364 266290 21416 266296
rect 18604 263560 18656 263566
rect 18604 263502 18656 263508
rect 18604 253972 18656 253978
rect 18604 253914 18656 253920
rect 18616 235958 18644 253914
rect 22744 252612 22796 252618
rect 22744 252554 22796 252560
rect 18604 235952 18656 235958
rect 18604 235894 18656 235900
rect 17224 215280 17276 215286
rect 17224 215222 17276 215228
rect 17224 186992 17276 186998
rect 17224 186934 17276 186940
rect 17236 111790 17264 186934
rect 17224 111784 17276 111790
rect 17224 111726 17276 111732
rect 22756 85542 22784 252554
rect 25516 150414 25544 289818
rect 29656 267714 29684 565830
rect 32416 287026 32444 670686
rect 39304 527196 39356 527202
rect 39304 527138 39356 527144
rect 33784 409896 33836 409902
rect 33784 409838 33836 409844
rect 32404 287020 32456 287026
rect 32404 286962 32456 286968
rect 32404 267776 32456 267782
rect 32404 267718 32456 267724
rect 29644 267708 29696 267714
rect 29644 267650 29696 267656
rect 25504 150408 25556 150414
rect 25504 150350 25556 150356
rect 22744 85536 22796 85542
rect 22744 85478 22796 85484
rect 23480 75200 23532 75206
rect 23480 75142 23532 75148
rect 19340 51740 19392 51746
rect 19340 51682 19392 51688
rect 15844 45552 15896 45558
rect 15844 45494 15896 45500
rect 16580 36576 16632 36582
rect 16580 36518 16632 36524
rect 16592 16574 16620 36518
rect 17960 19984 18012 19990
rect 17960 19926 18012 19932
rect 12452 16546 13584 16574
rect 13832 16546 14320 16574
rect 15212 16546 15976 16574
rect 16592 16546 17080 16574
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 11164 480 11192 15846
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11992 354 12020 3470
rect 13556 480 13584 16546
rect 12318 354 12430 480
rect 11992 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 15948 480 15976 16546
rect 17052 480 17080 16546
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 19926
rect 19352 16574 19380 51682
rect 20720 26920 20772 26926
rect 20720 26862 20772 26868
rect 20732 16574 20760 26862
rect 23492 16574 23520 75142
rect 30380 65544 30432 65550
rect 30380 65486 30432 65492
rect 29000 64184 29052 64190
rect 29000 64126 29052 64132
rect 27620 53100 27672 53106
rect 27620 53042 27672 53048
rect 24860 37936 24912 37942
rect 24860 37878 24912 37884
rect 24872 16574 24900 37878
rect 26240 28280 26292 28286
rect 26240 28222 26292 28228
rect 19352 16546 19472 16574
rect 20732 16546 21864 16574
rect 23492 16546 24256 16574
rect 24872 16546 25360 16574
rect 19444 480 19472 16546
rect 20168 14476 20220 14482
rect 20168 14418 20220 14424
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20180 354 20208 14418
rect 21836 480 21864 16546
rect 23020 3460 23072 3466
rect 23020 3402 23072 3408
rect 23032 480 23060 3402
rect 24228 480 24256 16546
rect 25332 480 25360 16546
rect 20598 354 20710 480
rect 20180 326 20710 354
rect 20598 -960 20710 326
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 28222
rect 27632 16574 27660 53042
rect 29012 16574 29040 64126
rect 30392 16574 30420 65486
rect 32416 33114 32444 267718
rect 33796 245614 33824 409838
rect 35164 397520 35216 397526
rect 35164 397462 35216 397468
rect 33784 245608 33836 245614
rect 33784 245550 33836 245556
rect 35176 237386 35204 397462
rect 39316 260846 39344 527138
rect 39304 260840 39356 260846
rect 39304 260782 39356 260788
rect 40052 238678 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 87604 703044 87656 703050
rect 87604 702986 87656 702992
rect 53748 702840 53800 702846
rect 53748 702782 53800 702788
rect 52368 590708 52420 590714
rect 52368 590650 52420 590656
rect 47584 462392 47636 462398
rect 47584 462334 47636 462340
rect 43444 371272 43496 371278
rect 43444 371214 43496 371220
rect 40040 238672 40092 238678
rect 40040 238614 40092 238620
rect 35164 237380 35216 237386
rect 35164 237322 35216 237328
rect 43456 235890 43484 371214
rect 47596 237318 47624 462334
rect 50344 294024 50396 294030
rect 50344 293966 50396 293972
rect 49608 270564 49660 270570
rect 49608 270506 49660 270512
rect 47584 237312 47636 237318
rect 47584 237254 47636 237260
rect 43444 235884 43496 235890
rect 43444 235826 43496 235832
rect 49620 210361 49648 270506
rect 49606 210352 49662 210361
rect 49606 210287 49662 210296
rect 50356 164218 50384 293966
rect 51724 278792 51776 278798
rect 51724 278734 51776 278740
rect 50988 257372 51040 257378
rect 50988 257314 51040 257320
rect 51000 211857 51028 257314
rect 50986 211848 51042 211857
rect 50986 211783 51042 211792
rect 50344 164212 50396 164218
rect 50344 164154 50396 164160
rect 44180 68332 44232 68338
rect 44180 68274 44232 68280
rect 34520 66904 34572 66910
rect 34520 66846 34572 66852
rect 33140 58676 33192 58682
rect 33140 58618 33192 58624
rect 32404 33108 32456 33114
rect 32404 33050 32456 33056
rect 31760 21412 31812 21418
rect 31760 21354 31812 21360
rect 31772 16574 31800 21354
rect 33152 16574 33180 58618
rect 27632 16546 28488 16574
rect 29012 16546 30144 16574
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 33152 16546 33640 16574
rect 27712 6180 27764 6186
rect 27712 6122 27764 6128
rect 27724 480 27752 6122
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28460 354 28488 16546
rect 30116 480 30144 16546
rect 28878 354 28990 480
rect 28460 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 33612 480 33640 16546
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 66846
rect 35898 62792 35954 62801
rect 35898 62727 35954 62736
rect 35912 3534 35940 62727
rect 35992 42084 36044 42090
rect 35992 42026 36044 42032
rect 35900 3528 35952 3534
rect 35900 3470 35952 3476
rect 36004 480 36032 42026
rect 42800 40724 42852 40730
rect 42800 40666 42852 40672
rect 40040 35284 40092 35290
rect 40040 35226 40092 35232
rect 37280 25560 37332 25566
rect 37280 25502 37332 25508
rect 37292 16574 37320 25502
rect 38660 17264 38712 17270
rect 38660 17206 38712 17212
rect 38672 16574 38700 17206
rect 40052 16574 40080 35226
rect 41420 24132 41472 24138
rect 41420 24074 41472 24080
rect 41432 16574 41460 24074
rect 37292 16546 38424 16574
rect 38672 16546 39160 16574
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 36820 3528 36872 3534
rect 36820 3470 36872 3476
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36832 354 36860 3470
rect 38396 480 38424 16546
rect 37158 354 37270 480
rect 36832 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 40666
rect 44192 3534 44220 68274
rect 45560 55956 45612 55962
rect 45560 55898 45612 55904
rect 44272 29640 44324 29646
rect 44272 29582 44324 29588
rect 44180 3528 44232 3534
rect 44180 3470 44232 3476
rect 44284 480 44312 29582
rect 45572 16574 45600 55898
rect 49698 47560 49754 47569
rect 49698 47495 49754 47504
rect 48320 33788 48372 33794
rect 48320 33730 48372 33736
rect 47582 32464 47638 32473
rect 47582 32399 47638 32408
rect 45572 16546 46704 16574
rect 45100 3528 45152 3534
rect 45100 3470 45152 3476
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45112 354 45140 3470
rect 46676 480 46704 16546
rect 47596 3466 47624 32399
rect 48332 16574 48360 33730
rect 49712 16574 49740 47495
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 47860 7608 47912 7614
rect 47860 7550 47912 7556
rect 47584 3460 47636 3466
rect 47584 3402 47636 3408
rect 47872 480 47900 7550
rect 45438 354 45550 480
rect 45112 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 51736 13190 51764 278734
rect 52380 238610 52408 590650
rect 53104 292800 53156 292806
rect 53104 292742 53156 292748
rect 52368 238604 52420 238610
rect 52368 238546 52420 238552
rect 53116 71738 53144 292742
rect 53656 264988 53708 264994
rect 53656 264930 53708 264936
rect 53668 217394 53696 264930
rect 53760 247042 53788 702782
rect 57888 702704 57940 702710
rect 57888 702646 57940 702652
rect 55128 700392 55180 700398
rect 55128 700334 55180 700340
rect 54484 357468 54536 357474
rect 54484 357410 54536 357416
rect 54496 312594 54524 357410
rect 54484 312588 54536 312594
rect 54484 312530 54536 312536
rect 54944 277432 54996 277438
rect 54944 277374 54996 277380
rect 53748 247036 53800 247042
rect 53748 246978 53800 246984
rect 54956 225622 54984 277374
rect 55036 276072 55088 276078
rect 55036 276014 55088 276020
rect 54944 225616 54996 225622
rect 54944 225558 54996 225564
rect 53656 217388 53708 217394
rect 53656 217330 53708 217336
rect 55048 188494 55076 276014
rect 55140 237250 55168 700334
rect 57796 282940 57848 282946
rect 57796 282882 57848 282888
rect 56416 277500 56468 277506
rect 56416 277442 56468 277448
rect 55128 237244 55180 237250
rect 55128 237186 55180 237192
rect 56428 207806 56456 277442
rect 57704 274712 57756 274718
rect 57704 274654 57756 274660
rect 56508 259480 56560 259486
rect 56508 259422 56560 259428
rect 56416 207800 56468 207806
rect 56416 207742 56468 207748
rect 55036 188488 55088 188494
rect 55036 188430 55088 188436
rect 56520 182850 56548 259422
rect 57520 258120 57572 258126
rect 57520 258062 57572 258068
rect 57532 194070 57560 258062
rect 57612 248464 57664 248470
rect 57612 248406 57664 248412
rect 57624 207738 57652 248406
rect 57612 207732 57664 207738
rect 57612 207674 57664 207680
rect 57716 199578 57744 274654
rect 57704 199572 57756 199578
rect 57704 199514 57756 199520
rect 57520 194064 57572 194070
rect 57520 194006 57572 194012
rect 57808 184278 57836 282882
rect 57900 255270 57928 702646
rect 62028 697672 62080 697678
rect 62028 697614 62080 697620
rect 59084 285728 59136 285734
rect 59084 285670 59136 285676
rect 57888 255264 57940 255270
rect 57888 255206 57940 255212
rect 58992 249824 59044 249830
rect 58992 249766 59044 249772
rect 59004 185638 59032 249766
rect 59096 218657 59124 285670
rect 61936 271992 61988 271998
rect 61936 271934 61988 271940
rect 60556 271924 60608 271930
rect 60556 271866 60608 271872
rect 59176 269136 59228 269142
rect 59176 269078 59228 269084
rect 59082 218648 59138 218657
rect 59082 218583 59138 218592
rect 59188 200802 59216 269078
rect 59268 263696 59320 263702
rect 59268 263638 59320 263644
rect 59176 200796 59228 200802
rect 59176 200738 59228 200744
rect 58992 185632 59044 185638
rect 58992 185574 59044 185580
rect 57796 184272 57848 184278
rect 57796 184214 57848 184220
rect 56508 182844 56560 182850
rect 56508 182786 56560 182792
rect 59280 180033 59308 263638
rect 60464 262268 60516 262274
rect 60464 262210 60516 262216
rect 60372 249892 60424 249898
rect 60372 249834 60424 249840
rect 60384 231266 60412 249834
rect 60372 231260 60424 231266
rect 60372 231202 60424 231208
rect 60476 213246 60504 262210
rect 60464 213240 60516 213246
rect 60464 213182 60516 213188
rect 60568 199510 60596 271866
rect 61844 260908 61896 260914
rect 61844 260850 61896 260856
rect 60648 255332 60700 255338
rect 60648 255274 60700 255280
rect 60556 199504 60608 199510
rect 60556 199446 60608 199452
rect 59266 180024 59322 180033
rect 59266 179959 59322 179968
rect 60660 178673 60688 255274
rect 61752 247104 61804 247110
rect 61752 247046 61804 247052
rect 61764 210458 61792 247046
rect 61856 221474 61884 260850
rect 61844 221468 61896 221474
rect 61844 221410 61896 221416
rect 61752 210452 61804 210458
rect 61752 210394 61804 210400
rect 61948 209098 61976 271934
rect 62040 249762 62068 697614
rect 66168 510672 66220 510678
rect 66168 510614 66220 510620
rect 63408 307828 63460 307834
rect 63408 307770 63460 307776
rect 63420 285666 63448 307770
rect 63408 285660 63460 285666
rect 63408 285602 63460 285608
rect 63408 280220 63460 280226
rect 63408 280162 63460 280168
rect 63316 251252 63368 251258
rect 63316 251194 63368 251200
rect 62028 249756 62080 249762
rect 62028 249698 62080 249704
rect 62028 247172 62080 247178
rect 62028 247114 62080 247120
rect 61936 209092 61988 209098
rect 61936 209034 61988 209040
rect 62040 191049 62068 247114
rect 63224 244316 63276 244322
rect 63224 244258 63276 244264
rect 63132 241528 63184 241534
rect 63132 241470 63184 241476
rect 63144 198014 63172 241470
rect 63236 233918 63264 244258
rect 63328 239494 63356 251194
rect 63316 239488 63368 239494
rect 63316 239430 63368 239436
rect 63224 233912 63276 233918
rect 63224 233854 63276 233860
rect 63420 204950 63448 280162
rect 66180 280158 66208 510614
rect 67548 404388 67600 404394
rect 67548 404330 67600 404336
rect 67456 294296 67508 294302
rect 67456 294238 67508 294244
rect 67468 291854 67496 294238
rect 67456 291848 67508 291854
rect 67456 291790 67508 291796
rect 67560 283121 67588 404330
rect 71792 308446 71820 702986
rect 79324 702500 79376 702506
rect 79324 702442 79376 702448
rect 75184 700324 75236 700330
rect 75184 700266 75236 700272
rect 75196 313993 75224 700266
rect 76564 351960 76616 351966
rect 76564 351902 76616 351908
rect 75182 313984 75238 313993
rect 75182 313919 75238 313928
rect 71780 308440 71832 308446
rect 71780 308382 71832 308388
rect 69020 305652 69072 305658
rect 69020 305594 69072 305600
rect 68650 300928 68706 300937
rect 68650 300863 68706 300872
rect 67638 290592 67694 290601
rect 67638 290527 67694 290536
rect 67652 289882 67680 290527
rect 67640 289876 67692 289882
rect 67640 289818 67692 289824
rect 68664 289785 68692 300863
rect 68834 296848 68890 296857
rect 68834 296783 68890 296792
rect 68744 295520 68796 295526
rect 68744 295462 68796 295468
rect 68756 290193 68784 295462
rect 68742 290184 68798 290193
rect 68742 290119 68798 290128
rect 68650 289776 68706 289785
rect 68650 289711 68706 289720
rect 68742 288824 68798 288833
rect 68742 288759 68798 288768
rect 67730 287056 67786 287065
rect 67640 287020 67692 287026
rect 67730 286991 67786 287000
rect 67640 286962 67692 286968
rect 67652 286793 67680 286962
rect 67638 286784 67694 286793
rect 67638 286719 67694 286728
rect 67744 285734 67772 286991
rect 68282 285832 68338 285841
rect 68282 285767 68338 285776
rect 67732 285728 67784 285734
rect 67732 285670 67784 285676
rect 67640 285660 67692 285666
rect 67640 285602 67692 285608
rect 67652 284753 67680 285602
rect 67638 284744 67694 284753
rect 67638 284679 67694 284688
rect 67638 283248 67694 283257
rect 67638 283183 67694 283192
rect 67546 283112 67602 283121
rect 67546 283047 67602 283056
rect 67652 282946 67680 283183
rect 67640 282940 67692 282946
rect 67640 282882 67692 282888
rect 67362 280528 67418 280537
rect 67362 280463 67418 280472
rect 66168 280152 66220 280158
rect 66168 280094 66220 280100
rect 65892 276140 65944 276146
rect 65892 276082 65944 276088
rect 63500 269816 63552 269822
rect 63500 269758 63552 269764
rect 63512 267646 63540 269758
rect 63500 267640 63552 267646
rect 63500 267582 63552 267588
rect 64788 258188 64840 258194
rect 64788 258130 64840 258136
rect 64604 255400 64656 255406
rect 64604 255342 64656 255348
rect 64512 245676 64564 245682
rect 64512 245618 64564 245624
rect 63500 239420 63552 239426
rect 63500 239362 63552 239368
rect 63512 238542 63540 239362
rect 63500 238536 63552 238542
rect 63500 238478 63552 238484
rect 63408 204944 63460 204950
rect 63408 204886 63460 204892
rect 63132 198008 63184 198014
rect 63132 197950 63184 197956
rect 64524 193866 64552 245618
rect 64616 203561 64644 255342
rect 64696 252680 64748 252686
rect 64696 252622 64748 252628
rect 64708 239562 64736 252622
rect 64696 239556 64748 239562
rect 64696 239498 64748 239504
rect 64602 203552 64658 203561
rect 64602 203487 64658 203496
rect 64512 193860 64564 193866
rect 64512 193802 64564 193808
rect 62026 191040 62082 191049
rect 62026 190975 62082 190984
rect 64800 188426 64828 258130
rect 64788 188420 64840 188426
rect 64788 188362 64840 188368
rect 65904 185774 65932 276082
rect 66076 273284 66128 273290
rect 66076 273226 66128 273232
rect 65984 260976 66036 260982
rect 65984 260918 66036 260924
rect 65996 194002 66024 260918
rect 66088 194138 66116 273226
rect 67270 269512 67326 269521
rect 67270 269447 67326 269456
rect 67284 228478 67312 269447
rect 67376 236706 67404 280463
rect 67638 280392 67694 280401
rect 67638 280327 67694 280336
rect 67652 280226 67680 280327
rect 67640 280220 67692 280226
rect 67640 280162 67692 280168
rect 67732 280152 67784 280158
rect 67732 280094 67784 280100
rect 67638 279168 67694 279177
rect 67638 279103 67694 279112
rect 67652 278798 67680 279103
rect 67744 279041 67772 280094
rect 67730 279032 67786 279041
rect 67730 278967 67786 278976
rect 67640 278792 67692 278798
rect 67640 278734 67692 278740
rect 67730 277808 67786 277817
rect 67730 277743 67786 277752
rect 67638 277672 67694 277681
rect 67638 277607 67694 277616
rect 67652 277506 67680 277607
rect 67640 277500 67692 277506
rect 67640 277442 67692 277448
rect 67744 277438 67772 277743
rect 67732 277432 67784 277438
rect 67732 277374 67784 277380
rect 67638 276448 67694 276457
rect 67638 276383 67694 276392
rect 67652 276078 67680 276383
rect 68006 276312 68062 276321
rect 68006 276247 68062 276256
rect 68020 276146 68048 276247
rect 68008 276140 68060 276146
rect 68008 276082 68060 276088
rect 67640 276072 67692 276078
rect 67640 276014 67692 276020
rect 67638 275088 67694 275097
rect 67638 275023 67694 275032
rect 67652 274718 67680 275023
rect 67640 274712 67692 274718
rect 67640 274654 67692 274660
rect 67732 274644 67784 274650
rect 67732 274586 67784 274592
rect 67744 274553 67772 274586
rect 67730 274544 67786 274553
rect 67730 274479 67786 274488
rect 68006 273592 68062 273601
rect 68006 273527 68062 273536
rect 68020 273290 68048 273527
rect 68008 273284 68060 273290
rect 68008 273226 68060 273232
rect 67730 272368 67786 272377
rect 67730 272303 67786 272312
rect 67638 272232 67694 272241
rect 67638 272167 67694 272176
rect 67652 271998 67680 272167
rect 67640 271992 67692 271998
rect 67640 271934 67692 271940
rect 67744 271930 67772 272303
rect 67732 271924 67784 271930
rect 67732 271866 67784 271872
rect 67638 271008 67694 271017
rect 67638 270943 67694 270952
rect 67652 270570 67680 270943
rect 67640 270564 67692 270570
rect 67640 270506 67692 270512
rect 67638 269648 67694 269657
rect 67638 269583 67694 269592
rect 67652 269142 67680 269583
rect 67640 269136 67692 269142
rect 67640 269078 67692 269084
rect 67638 268152 67694 268161
rect 67638 268087 67694 268096
rect 67652 267782 67680 268087
rect 67640 267776 67692 267782
rect 67640 267718 67692 267724
rect 67732 267708 67784 267714
rect 67732 267650 67784 267656
rect 67640 267640 67692 267646
rect 67640 267582 67692 267588
rect 67652 267073 67680 267582
rect 67744 267481 67772 267650
rect 67730 267472 67786 267481
rect 67730 267407 67786 267416
rect 67638 267064 67694 267073
rect 67638 266999 67694 267008
rect 67732 266348 67784 266354
rect 67732 266290 67784 266296
rect 67638 265432 67694 265441
rect 67638 265367 67694 265376
rect 67652 264994 67680 265367
rect 67744 265033 67772 266290
rect 67730 265024 67786 265033
rect 67640 264988 67692 264994
rect 67730 264959 67786 264968
rect 67640 264930 67692 264936
rect 67730 264208 67786 264217
rect 67730 264143 67786 264152
rect 67640 263696 67692 263702
rect 67638 263664 67640 263673
rect 67692 263664 67694 263673
rect 67744 263634 67772 264143
rect 67638 263599 67694 263608
rect 67732 263628 67784 263634
rect 67732 263570 67784 263576
rect 67640 263560 67692 263566
rect 67638 263528 67640 263537
rect 67692 263528 67694 263537
rect 67638 263463 67694 263472
rect 67638 262304 67694 262313
rect 67638 262239 67640 262248
rect 67692 262239 67694 262248
rect 67640 262210 67692 262216
rect 67730 261488 67786 261497
rect 67730 261423 67786 261432
rect 67640 260976 67692 260982
rect 67638 260944 67640 260953
rect 67692 260944 67694 260953
rect 67744 260914 67772 261423
rect 67638 260879 67694 260888
rect 67732 260908 67784 260914
rect 67732 260850 67784 260856
rect 67640 260840 67692 260846
rect 67638 260808 67640 260817
rect 67692 260808 67694 260817
rect 67638 260743 67694 260752
rect 67638 259584 67694 259593
rect 67638 259519 67694 259528
rect 67652 259486 67680 259519
rect 67640 259480 67692 259486
rect 67640 259422 67692 259428
rect 67730 258632 67786 258641
rect 67730 258567 67786 258576
rect 67638 258224 67694 258233
rect 67638 258159 67640 258168
rect 67692 258159 67694 258168
rect 67640 258130 67692 258136
rect 67744 258126 67772 258567
rect 67732 258120 67784 258126
rect 67732 258062 67784 258068
rect 68296 257378 68324 285767
rect 68756 282169 68784 288759
rect 68848 288153 68876 296783
rect 68928 292596 68980 292602
rect 68928 292538 68980 292544
rect 68940 289513 68968 292538
rect 68926 289504 68982 289513
rect 68926 289439 68982 289448
rect 68834 288144 68890 288153
rect 68834 288079 68890 288088
rect 68742 282160 68798 282169
rect 68742 282095 68798 282104
rect 68374 275224 68430 275233
rect 68374 275159 68430 275168
rect 68284 257372 68336 257378
rect 68284 257314 68336 257320
rect 67638 257272 67694 257281
rect 67638 257207 67694 257216
rect 67652 256766 67680 257207
rect 67640 256760 67692 256766
rect 67640 256702 67692 256708
rect 67638 255912 67694 255921
rect 67638 255847 67694 255856
rect 67652 255406 67680 255847
rect 67640 255400 67692 255406
rect 67640 255342 67692 255348
rect 67730 255368 67786 255377
rect 67730 255303 67732 255312
rect 67784 255303 67786 255312
rect 67732 255274 67784 255280
rect 67640 255264 67692 255270
rect 67638 255232 67640 255241
rect 67692 255232 67694 255241
rect 67638 255167 67694 255176
rect 67730 253192 67786 253201
rect 67730 253127 67786 253136
rect 67638 252784 67694 252793
rect 67638 252719 67694 252728
rect 67652 252686 67680 252719
rect 67640 252680 67692 252686
rect 67640 252622 67692 252628
rect 67744 252618 67772 253127
rect 67732 252612 67784 252618
rect 67732 252554 67784 252560
rect 67638 251832 67694 251841
rect 67638 251767 67694 251776
rect 67652 251258 67680 251767
rect 67640 251252 67692 251258
rect 67640 251194 67692 251200
rect 67730 250472 67786 250481
rect 67730 250407 67786 250416
rect 67638 249928 67694 249937
rect 67638 249863 67640 249872
rect 67692 249863 67694 249872
rect 67640 249834 67692 249840
rect 67744 249830 67772 250407
rect 67732 249824 67784 249830
rect 67638 249792 67694 249801
rect 67732 249766 67784 249772
rect 67638 249727 67640 249736
rect 67692 249727 67694 249736
rect 67640 249698 67692 249704
rect 68388 249694 68416 275159
rect 69032 270881 69060 305594
rect 70400 305040 70452 305046
rect 70400 304982 70452 304988
rect 75920 305040 75972 305046
rect 75920 304982 75972 304988
rect 69664 302388 69716 302394
rect 69664 302330 69716 302336
rect 69676 291938 69704 302330
rect 70412 301510 70440 304982
rect 74540 303680 74592 303686
rect 74540 303622 74592 303628
rect 71780 302252 71832 302258
rect 71780 302194 71832 302200
rect 70400 301504 70452 301510
rect 70400 301446 70452 301452
rect 70400 301368 70452 301374
rect 70400 301310 70452 301316
rect 70412 294370 70440 301310
rect 70492 299600 70544 299606
rect 70492 299542 70544 299548
rect 70400 294364 70452 294370
rect 70400 294306 70452 294312
rect 70504 291977 70532 299542
rect 71044 294364 71096 294370
rect 71044 294306 71096 294312
rect 71056 291977 71084 294306
rect 71792 291977 71820 302194
rect 72608 298784 72660 298790
rect 72608 298726 72660 298732
rect 70504 291949 70702 291977
rect 71056 291949 71346 291977
rect 71792 291949 71990 291977
rect 72620 291963 72648 298726
rect 73896 298172 73948 298178
rect 73896 298114 73948 298120
rect 73252 294636 73304 294642
rect 73252 294578 73304 294584
rect 73264 291963 73292 294578
rect 73908 291963 73936 298114
rect 74552 291963 74580 303622
rect 75184 295452 75236 295458
rect 75184 295394 75236 295400
rect 75196 291963 75224 295394
rect 75826 294264 75882 294273
rect 75826 294199 75882 294208
rect 75840 291963 75868 294199
rect 75932 291977 75960 304982
rect 76576 298178 76604 351902
rect 77300 313948 77352 313954
rect 77300 313890 77352 313896
rect 77312 306374 77340 313890
rect 77312 306346 78076 306374
rect 76564 298172 76616 298178
rect 76564 298114 76616 298120
rect 77116 296744 77168 296750
rect 77116 296686 77168 296692
rect 75932 291949 76498 291977
rect 77128 291963 77156 296686
rect 77760 294364 77812 294370
rect 77760 294306 77812 294312
rect 77772 291963 77800 294306
rect 78048 291938 78076 306346
rect 79336 294370 79364 702442
rect 84476 304292 84528 304298
rect 84476 304234 84528 304240
rect 81900 303748 81952 303754
rect 81900 303690 81952 303696
rect 80060 299532 80112 299538
rect 80060 299474 80112 299480
rect 79692 298376 79744 298382
rect 79692 298318 79744 298324
rect 79324 294364 79376 294370
rect 79324 294306 79376 294312
rect 79048 294024 79100 294030
rect 79048 293966 79100 293972
rect 79060 291963 79088 293966
rect 79704 291963 79732 298318
rect 80072 291977 80100 299474
rect 81624 294024 81676 294030
rect 81624 293966 81676 293972
rect 80980 292664 81032 292670
rect 80980 292606 81032 292612
rect 80072 291949 80362 291977
rect 80992 291963 81020 292606
rect 81636 291963 81664 293966
rect 81912 291938 81940 303690
rect 84292 299668 84344 299674
rect 84292 299610 84344 299616
rect 83556 298308 83608 298314
rect 83556 298250 83608 298256
rect 82912 297016 82964 297022
rect 82912 296958 82964 296964
rect 82924 291963 82952 296958
rect 83568 291963 83596 298250
rect 84304 291977 84332 299610
rect 84226 291949 84332 291977
rect 84488 291938 84516 304234
rect 85580 303816 85632 303822
rect 85580 303758 85632 303764
rect 85488 295112 85540 295118
rect 85488 295054 85540 295060
rect 85500 291963 85528 295054
rect 85592 294370 85620 303758
rect 85672 300960 85724 300966
rect 85672 300902 85724 300908
rect 85580 294364 85632 294370
rect 85580 294306 85632 294312
rect 85684 291938 85712 300902
rect 87616 295118 87644 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 88352 327758 88380 702406
rect 105464 700398 105492 703520
rect 107660 702976 107712 702982
rect 107660 702918 107712 702924
rect 106280 702772 106332 702778
rect 106280 702714 106332 702720
rect 105452 700392 105504 700398
rect 105452 700334 105504 700340
rect 97264 563100 97316 563106
rect 97264 563042 97316 563048
rect 93124 418192 93176 418198
rect 93124 418134 93176 418140
rect 88340 327752 88392 327758
rect 88340 327694 88392 327700
rect 91100 319456 91152 319462
rect 91100 319398 91152 319404
rect 89720 306400 89772 306406
rect 89720 306342 89772 306348
rect 89352 298512 89404 298518
rect 89352 298454 89404 298460
rect 88708 298172 88760 298178
rect 88708 298114 88760 298120
rect 88064 295588 88116 295594
rect 88064 295530 88116 295536
rect 87604 295112 87656 295118
rect 87604 295054 87656 295060
rect 86500 294364 86552 294370
rect 86500 294306 86552 294312
rect 86512 291977 86540 294306
rect 87420 294228 87472 294234
rect 87420 294170 87472 294176
rect 86512 291949 86802 291977
rect 87432 291963 87460 294170
rect 88076 291963 88104 295530
rect 88720 291963 88748 298114
rect 89364 291963 89392 298454
rect 89732 291977 89760 306342
rect 90364 302456 90416 302462
rect 90364 302398 90416 302404
rect 90376 291977 90404 302398
rect 91112 291977 91140 319398
rect 93136 313954 93164 418134
rect 97276 317558 97304 563042
rect 101404 345092 101456 345098
rect 101404 345034 101456 345040
rect 93952 317552 94004 317558
rect 93952 317494 94004 317500
rect 97264 317552 97316 317558
rect 97264 317494 97316 317500
rect 93124 313948 93176 313954
rect 93124 313890 93176 313896
rect 92664 305108 92716 305114
rect 92664 305050 92716 305056
rect 92572 294296 92624 294302
rect 92572 294238 92624 294244
rect 91928 294160 91980 294166
rect 91928 294102 91980 294108
rect 89732 291949 90022 291977
rect 90376 291949 90666 291977
rect 91112 291949 91310 291977
rect 91940 291963 91968 294102
rect 92584 291963 92612 294238
rect 92676 291977 92704 305050
rect 93964 294370 93992 317494
rect 98000 312588 98052 312594
rect 98000 312530 98052 312536
rect 94136 311160 94188 311166
rect 94136 311102 94188 311108
rect 93952 294364 94004 294370
rect 93952 294306 94004 294312
rect 93860 292732 93912 292738
rect 93860 292674 93912 292680
rect 92676 291949 93242 291977
rect 93872 291963 93900 292674
rect 94148 291977 94176 311102
rect 97724 296812 97776 296818
rect 97724 296754 97776 296760
rect 94780 294364 94832 294370
rect 94780 294306 94832 294312
rect 94148 291949 94530 291977
rect 94792 291938 94820 294306
rect 95790 294128 95846 294137
rect 95790 294063 95846 294072
rect 97080 294092 97132 294098
rect 95804 291963 95832 294063
rect 97080 294034 97132 294040
rect 96436 292868 96488 292874
rect 96436 292810 96488 292816
rect 96448 291963 96476 292810
rect 97092 291963 97120 294034
rect 97736 291963 97764 296754
rect 98012 291977 98040 312530
rect 101416 311166 101444 345034
rect 103796 327752 103848 327758
rect 103796 327694 103848 327700
rect 101404 311160 101456 311166
rect 101404 311102 101456 311108
rect 103808 306374 103836 327694
rect 106292 306374 106320 702714
rect 107672 306374 107700 702918
rect 129004 702908 129056 702914
rect 129004 702850 129056 702856
rect 124864 702636 124916 702642
rect 124864 702578 124916 702584
rect 123484 643136 123536 643142
rect 123484 643078 123536 643084
rect 116584 579692 116636 579698
rect 116584 579634 116636 579640
rect 111064 474768 111116 474774
rect 111064 474710 111116 474716
rect 103808 306346 104296 306374
rect 106292 306346 106872 306374
rect 107672 306346 108344 306374
rect 100852 302320 100904 302326
rect 100852 302262 100904 302268
rect 99656 295724 99708 295730
rect 99656 295666 99708 295672
rect 99012 295384 99064 295390
rect 99012 295326 99064 295332
rect 98012 291949 98394 291977
rect 99024 291963 99052 295326
rect 99668 291963 99696 295666
rect 100864 291977 100892 302262
rect 102140 300892 102192 300898
rect 102140 300834 102192 300840
rect 101588 292800 101640 292806
rect 101588 292742 101640 292748
rect 100864 291949 100970 291977
rect 101600 291963 101628 292742
rect 102152 291977 102180 300834
rect 102324 299736 102376 299742
rect 102324 299678 102376 299684
rect 102152 291949 102258 291977
rect 102336 291938 102364 299678
rect 103520 292800 103572 292806
rect 103520 292742 103572 292748
rect 103532 291963 103560 292742
rect 104162 292632 104218 292641
rect 104162 292567 104218 292576
rect 104176 291963 104204 292567
rect 104268 291977 104296 306346
rect 106094 298208 106150 298217
rect 106094 298143 106150 298152
rect 105450 292768 105506 292777
rect 105450 292703 105506 292712
rect 104268 291949 104834 291977
rect 105464 291963 105492 292703
rect 106108 291963 106136 298143
rect 106740 294364 106792 294370
rect 106740 294306 106792 294312
rect 106752 291963 106780 294306
rect 106844 291977 106872 306346
rect 108316 291977 108344 306346
rect 110604 298444 110656 298450
rect 110604 298386 110656 298392
rect 109958 295352 110014 295361
rect 109958 295287 110014 295296
rect 109316 292868 109368 292874
rect 109316 292810 109368 292816
rect 106844 291949 107410 291977
rect 108210 291952 108266 291961
rect 69676 291910 70058 291938
rect 78048 291910 78418 291938
rect 81912 291910 82282 291938
rect 84488 291910 84858 291938
rect 85684 291910 86146 291938
rect 94792 291910 95162 291938
rect 102336 291910 102890 291938
rect 108054 291910 108210 291938
rect 108316 291949 108698 291977
rect 109328 291963 109356 292810
rect 109972 291963 110000 295287
rect 110616 291963 110644 298386
rect 111076 293282 111104 474710
rect 116596 318782 116624 579634
rect 120080 501016 120132 501022
rect 120080 500958 120132 500964
rect 116584 318776 116636 318782
rect 116584 318718 116636 318724
rect 115940 318096 115992 318102
rect 115940 318038 115992 318044
rect 114560 308440 114612 308446
rect 114560 308382 114612 308388
rect 111248 298240 111300 298246
rect 111248 298182 111300 298188
rect 111064 293276 111116 293282
rect 111064 293218 111116 293224
rect 111260 291963 111288 298182
rect 112536 297084 112588 297090
rect 112536 297026 112588 297032
rect 111798 295488 111854 295497
rect 111798 295423 111854 295432
rect 111812 294642 111840 295423
rect 111800 294636 111852 294642
rect 111800 294578 111852 294584
rect 111892 294296 111944 294302
rect 111892 294238 111944 294244
rect 111904 291963 111932 294238
rect 112548 291963 112576 297026
rect 113824 296880 113876 296886
rect 113824 296822 113876 296828
rect 113178 293992 113234 294001
rect 113178 293927 113234 293936
rect 113192 291963 113220 293927
rect 113836 291963 113864 296822
rect 114468 294092 114520 294098
rect 114468 294034 114520 294040
rect 114480 291963 114508 294034
rect 114572 291977 114600 308382
rect 115952 291977 115980 318038
rect 118700 311160 118752 311166
rect 118700 311102 118752 311108
rect 118712 306374 118740 311102
rect 118712 306346 119200 306374
rect 117688 296948 117740 296954
rect 117688 296890 117740 296896
rect 114572 291949 115138 291977
rect 115952 291949 116426 291977
rect 117700 291963 117728 296890
rect 118332 295656 118384 295662
rect 118332 295598 118384 295604
rect 118344 291963 118372 295598
rect 119068 291984 119120 291990
rect 119002 291949 119068 291977
rect 117070 291922 117268 291938
rect 119068 291926 119120 291932
rect 119172 291938 119200 306346
rect 119712 294364 119764 294370
rect 119712 294306 119764 294312
rect 108210 291887 108266 291896
rect 115848 291916 115900 291922
rect 115782 291864 115848 291870
rect 117070 291916 117280 291922
rect 117070 291910 117228 291916
rect 115782 291858 115900 291864
rect 119172 291910 119646 291938
rect 117228 291858 117280 291864
rect 115782 291842 115888 291858
rect 69754 291272 69810 291281
rect 69754 291207 69756 291216
rect 69808 291207 69810 291216
rect 69756 291178 69808 291184
rect 119724 287054 119752 294306
rect 119804 291984 119856 291990
rect 119804 291926 119856 291932
rect 119816 290601 119844 291926
rect 119802 290592 119858 290601
rect 119802 290527 119858 290536
rect 119724 287026 119844 287054
rect 69018 270872 69074 270881
rect 69018 270807 69074 270816
rect 69202 268288 69258 268297
rect 69202 268223 69258 268232
rect 69110 251288 69166 251297
rect 69110 251223 69166 251232
rect 67548 249688 67600 249694
rect 67548 249630 67600 249636
rect 68376 249688 68428 249694
rect 68376 249630 68428 249636
rect 67454 240272 67510 240281
rect 67454 240207 67510 240216
rect 67364 236700 67416 236706
rect 67364 236642 67416 236648
rect 67272 228472 67324 228478
rect 67272 228414 67324 228420
rect 66076 194132 66128 194138
rect 66076 194074 66128 194080
rect 65984 193996 66036 194002
rect 65984 193938 66036 193944
rect 65892 185768 65944 185774
rect 65892 185710 65944 185716
rect 67468 180130 67496 240207
rect 67560 185706 67588 249630
rect 67638 248568 67694 248577
rect 67638 248503 67694 248512
rect 67652 248470 67680 248503
rect 67640 248464 67692 248470
rect 67640 248406 67692 248412
rect 67638 247752 67694 247761
rect 67638 247687 67694 247696
rect 67652 247178 67680 247687
rect 67730 247208 67786 247217
rect 67640 247172 67692 247178
rect 67730 247143 67786 247152
rect 67640 247114 67692 247120
rect 67744 247110 67772 247143
rect 67732 247104 67784 247110
rect 67732 247046 67784 247052
rect 67640 247036 67692 247042
rect 67640 246978 67692 246984
rect 67652 246673 67680 246978
rect 67638 246664 67694 246673
rect 67638 246599 67694 246608
rect 67730 245984 67786 245993
rect 67730 245919 67786 245928
rect 67744 245682 67772 245919
rect 67732 245676 67784 245682
rect 67732 245618 67784 245624
rect 67640 245608 67692 245614
rect 67640 245550 67692 245556
rect 67652 245313 67680 245550
rect 67638 245304 67694 245313
rect 67638 245239 67694 245248
rect 67638 244624 67694 244633
rect 67638 244559 67694 244568
rect 67652 244322 67680 244559
rect 67640 244316 67692 244322
rect 67640 244258 67692 244264
rect 67732 244248 67784 244254
rect 67732 244190 67784 244196
rect 67744 243953 67772 244190
rect 67730 243944 67786 243953
rect 67730 243879 67786 243888
rect 67638 241904 67694 241913
rect 67638 241839 67694 241848
rect 67652 241534 67680 241839
rect 67640 241528 67692 241534
rect 67640 241470 67692 241476
rect 69020 233980 69072 233986
rect 69020 233922 69072 233928
rect 67548 185700 67600 185706
rect 67548 185642 67600 185648
rect 69032 184210 69060 233922
rect 69124 196625 69152 251223
rect 69216 232558 69244 268223
rect 119816 261526 119844 287026
rect 120092 268705 120120 500958
rect 120264 324964 120316 324970
rect 120264 324906 120316 324912
rect 120172 315308 120224 315314
rect 120172 315250 120224 315256
rect 120078 268696 120134 268705
rect 120078 268631 120134 268640
rect 119804 261520 119856 261526
rect 119804 261462 119856 261468
rect 120078 251016 120134 251025
rect 120078 250951 120134 250960
rect 69662 244216 69718 244225
rect 69662 244151 69718 244160
rect 69676 239426 69704 244151
rect 119802 240952 119858 240961
rect 119802 240887 119858 240896
rect 69768 240094 70058 240122
rect 119646 240094 119752 240122
rect 69664 239420 69716 239426
rect 69664 239362 69716 239368
rect 69768 233986 69796 240094
rect 70688 238754 70716 240037
rect 70412 238726 70716 238754
rect 69756 233980 69808 233986
rect 69756 233922 69808 233928
rect 69204 232552 69256 232558
rect 69204 232494 69256 232500
rect 69110 196616 69166 196625
rect 69110 196551 69166 196560
rect 70412 188358 70440 238726
rect 71332 238066 71360 240037
rect 71976 238754 72004 240037
rect 72424 239556 72476 239562
rect 72424 239498 72476 239504
rect 71792 238726 72004 238754
rect 71320 238060 71372 238066
rect 71320 238002 71372 238008
rect 70400 188352 70452 188358
rect 70400 188294 70452 188300
rect 69020 184204 69072 184210
rect 69020 184146 69072 184152
rect 71792 182889 71820 238726
rect 71778 182880 71834 182889
rect 71778 182815 71834 182824
rect 72436 180198 72464 239498
rect 72620 238134 72648 240037
rect 73160 239828 73212 239834
rect 73160 239770 73212 239776
rect 72608 238128 72660 238134
rect 72608 238070 72660 238076
rect 73172 189786 73200 239770
rect 73264 225593 73292 240037
rect 73896 239834 73924 240037
rect 73884 239828 73936 239834
rect 73884 239770 73936 239776
rect 74552 238754 74580 240037
rect 75196 238754 75224 240037
rect 74552 238726 74672 238754
rect 73250 225584 73306 225593
rect 73250 225519 73306 225528
rect 74644 214606 74672 238726
rect 74736 238726 75224 238754
rect 74632 214600 74684 214606
rect 74632 214542 74684 214548
rect 73160 189780 73212 189786
rect 73160 189722 73212 189728
rect 74736 181490 74764 238726
rect 75840 238610 75868 240037
rect 75920 239828 75972 239834
rect 75920 239770 75972 239776
rect 75828 238604 75880 238610
rect 75828 238546 75880 238552
rect 75932 217326 75960 239770
rect 76484 238754 76512 240037
rect 77116 239834 77144 240037
rect 77104 239828 77156 239834
rect 77104 239770 77156 239776
rect 77300 239828 77352 239834
rect 77300 239770 77352 239776
rect 76024 238726 76512 238754
rect 76024 228410 76052 238726
rect 76012 228404 76064 228410
rect 76012 228346 76064 228352
rect 75920 217320 75972 217326
rect 75920 217262 75972 217268
rect 77312 206378 77340 239770
rect 77772 238754 77800 240037
rect 78404 239834 78432 240037
rect 78392 239828 78444 239834
rect 78392 239770 78444 239776
rect 78680 239828 78732 239834
rect 78680 239770 78732 239776
rect 77404 238726 77800 238754
rect 77404 218754 77432 238726
rect 77392 218748 77444 218754
rect 77392 218690 77444 218696
rect 78692 207670 78720 239770
rect 79060 238754 79088 240037
rect 79692 239834 79720 240037
rect 79680 239828 79732 239834
rect 79680 239770 79732 239776
rect 78784 238726 79088 238754
rect 78784 216034 78812 238726
rect 79324 238060 79376 238066
rect 79324 238002 79376 238008
rect 78772 216028 78824 216034
rect 78772 215970 78824 215976
rect 78680 207664 78732 207670
rect 78680 207606 78732 207612
rect 77300 206372 77352 206378
rect 77300 206314 77352 206320
rect 79336 192545 79364 238002
rect 80348 235346 80376 240037
rect 80980 239816 81008 240037
rect 80900 239788 81008 239816
rect 80336 235340 80388 235346
rect 80336 235282 80388 235288
rect 80900 219434 80928 239788
rect 81636 238202 81664 240037
rect 81624 238196 81676 238202
rect 81624 238138 81676 238144
rect 82280 237386 82308 240037
rect 82820 239828 82872 239834
rect 82820 239770 82872 239776
rect 82268 237380 82320 237386
rect 82268 237322 82320 237328
rect 80072 219406 80928 219434
rect 79322 192536 79378 192545
rect 79322 192471 79378 192480
rect 80072 185842 80100 219406
rect 80060 185836 80112 185842
rect 80060 185778 80112 185784
rect 74724 181484 74776 181490
rect 74724 181426 74776 181432
rect 72424 180192 72476 180198
rect 72424 180134 72476 180140
rect 67456 180124 67508 180130
rect 67456 180066 67508 180072
rect 60646 178664 60702 178673
rect 60646 178599 60702 178608
rect 82832 177342 82860 239770
rect 82924 224330 82952 240037
rect 83556 239834 83584 240037
rect 83544 239828 83596 239834
rect 83544 239770 83596 239776
rect 84212 239442 84240 240037
rect 84212 239414 84424 239442
rect 84292 239352 84344 239358
rect 84292 239294 84344 239300
rect 84108 231872 84160 231878
rect 84160 231826 84240 231854
rect 84108 231814 84160 231820
rect 82912 224324 82964 224330
rect 82912 224266 82964 224272
rect 84212 191350 84240 231826
rect 84304 222902 84332 239294
rect 84292 222896 84344 222902
rect 84396 222873 84424 239414
rect 84856 231878 84884 240037
rect 85500 239358 85528 240037
rect 85488 239352 85540 239358
rect 85488 239294 85540 239300
rect 86144 238066 86172 240037
rect 86788 238542 86816 240037
rect 86960 239828 87012 239834
rect 86960 239770 87012 239776
rect 86776 238536 86828 238542
rect 86776 238478 86828 238484
rect 86132 238060 86184 238066
rect 86132 238002 86184 238008
rect 84844 231872 84896 231878
rect 84844 231814 84896 231820
rect 84292 222838 84344 222844
rect 84382 222864 84438 222873
rect 84382 222799 84438 222808
rect 86972 195362 87000 239770
rect 87432 238754 87460 240037
rect 88064 239834 88092 240037
rect 88052 239828 88104 239834
rect 88052 239770 88104 239776
rect 88720 238754 88748 240037
rect 87064 238726 87460 238754
rect 88444 238726 88748 238754
rect 87064 199442 87092 238726
rect 87052 199436 87104 199442
rect 87052 199378 87104 199384
rect 86960 195356 87012 195362
rect 86960 195298 87012 195304
rect 88444 193934 88472 238726
rect 89364 237250 89392 240037
rect 89720 239828 89772 239834
rect 89720 239770 89772 239776
rect 89352 237244 89404 237250
rect 89352 237186 89404 237192
rect 89732 198082 89760 239770
rect 90008 238754 90036 240037
rect 90640 239834 90668 240037
rect 90628 239828 90680 239834
rect 90628 239770 90680 239776
rect 89824 238726 90036 238754
rect 89824 221542 89852 238726
rect 91296 238610 91324 240037
rect 91284 238604 91336 238610
rect 91284 238546 91336 238552
rect 91100 238128 91152 238134
rect 91100 238070 91152 238076
rect 91112 230450 91140 238070
rect 91940 234598 91968 240037
rect 92480 239828 92532 239834
rect 92480 239770 92532 239776
rect 91928 234592 91980 234598
rect 91928 234534 91980 234540
rect 91100 230444 91152 230450
rect 91100 230386 91152 230392
rect 89812 221536 89864 221542
rect 89812 221478 89864 221484
rect 89720 198076 89772 198082
rect 89720 198018 89772 198024
rect 88432 193928 88484 193934
rect 88432 193870 88484 193876
rect 84200 191344 84252 191350
rect 84200 191286 84252 191292
rect 92492 188329 92520 239770
rect 92584 191418 92612 240037
rect 93216 239834 93244 240037
rect 93204 239828 93256 239834
rect 93204 239770 93256 239776
rect 93872 233866 93900 240037
rect 94516 238754 94544 240037
rect 95148 239850 95176 240037
rect 94056 238726 94544 238754
rect 95068 239822 95176 239850
rect 93872 233838 93992 233866
rect 93860 233776 93912 233782
rect 93860 233718 93912 233724
rect 92572 191412 92624 191418
rect 92572 191354 92624 191360
rect 92478 188320 92534 188329
rect 92478 188255 92534 188264
rect 93872 182918 93900 233718
rect 93964 209166 93992 233838
rect 94056 233782 94084 238726
rect 94044 233776 94096 233782
rect 94044 233718 94096 233724
rect 95068 219434 95096 239822
rect 95804 238678 95832 240037
rect 96436 239850 96464 240037
rect 96356 239822 96464 239850
rect 95792 238672 95844 238678
rect 95792 238614 95844 238620
rect 96356 219434 96384 239822
rect 97092 238754 97120 240037
rect 97724 239850 97752 240037
rect 94056 219406 95096 219434
rect 95344 219406 96384 219434
rect 96632 238726 97120 238754
rect 97644 239822 97752 239850
rect 94056 215966 94084 219406
rect 94044 215960 94096 215966
rect 94044 215902 94096 215908
rect 93952 209160 94004 209166
rect 93952 209102 94004 209108
rect 95344 191214 95372 219406
rect 96632 211818 96660 238726
rect 97644 224262 97672 239822
rect 98380 237386 98408 240037
rect 98644 239488 98696 239494
rect 98644 239430 98696 239436
rect 98368 237380 98420 237386
rect 98368 237322 98420 237328
rect 97632 224256 97684 224262
rect 97632 224198 97684 224204
rect 96620 211812 96672 211818
rect 96620 211754 96672 211760
rect 98656 206310 98684 239430
rect 99024 235890 99052 240037
rect 99668 238754 99696 240037
rect 100300 239850 100328 240037
rect 99392 238726 99696 238754
rect 100220 239822 100328 239850
rect 99012 235884 99064 235890
rect 99012 235826 99064 235832
rect 98644 206304 98696 206310
rect 98644 206246 98696 206252
rect 99392 195294 99420 238726
rect 100220 219434 100248 239822
rect 100956 238754 100984 240037
rect 101588 239850 101616 240037
rect 102232 239850 102260 240037
rect 99484 219406 100248 219434
rect 100772 238726 100984 238754
rect 101508 239822 101616 239850
rect 102152 239822 102260 239850
rect 99484 196654 99512 219406
rect 100772 203658 100800 238726
rect 101508 219434 101536 239822
rect 100864 219406 101536 219434
rect 100864 214674 100892 219406
rect 100852 214668 100904 214674
rect 100852 214610 100904 214616
rect 100760 203652 100812 203658
rect 100760 203594 100812 203600
rect 99472 196648 99524 196654
rect 99472 196590 99524 196596
rect 99380 195288 99432 195294
rect 99380 195230 99432 195236
rect 95332 191208 95384 191214
rect 95332 191150 95384 191156
rect 102152 191146 102180 239822
rect 102888 238270 102916 240037
rect 103532 238746 103560 240037
rect 104176 238754 104204 240037
rect 104808 239850 104836 240037
rect 103520 238740 103572 238746
rect 103520 238682 103572 238688
rect 103624 238726 104204 238754
rect 104728 239822 104836 239850
rect 104900 239828 104952 239834
rect 102876 238264 102928 238270
rect 102876 238206 102928 238212
rect 103624 205086 103652 238726
rect 104728 219434 104756 239822
rect 104900 239770 104952 239776
rect 103716 219406 104756 219434
rect 103612 205080 103664 205086
rect 103612 205022 103664 205028
rect 103716 202230 103744 219406
rect 103704 202224 103756 202230
rect 103704 202166 103756 202172
rect 104912 202162 104940 239770
rect 105464 238134 105492 240037
rect 106096 239834 106124 240037
rect 106084 239828 106136 239834
rect 106084 239770 106136 239776
rect 106752 238814 106780 240037
rect 106740 238808 106792 238814
rect 106740 238750 106792 238756
rect 107396 238754 107424 240037
rect 108040 238754 108068 240037
rect 108672 239850 108700 240037
rect 109960 239850 109988 240037
rect 106844 238726 107424 238754
rect 107672 238726 108068 238754
rect 108592 239822 108700 239850
rect 109880 239822 109988 239850
rect 105452 238128 105504 238134
rect 105452 238070 105504 238076
rect 106844 231810 106872 238726
rect 106924 238264 106976 238270
rect 106924 238206 106976 238212
rect 106832 231804 106884 231810
rect 106832 231746 106884 231752
rect 104900 202156 104952 202162
rect 104900 202098 104952 202104
rect 106936 192506 106964 238206
rect 106924 192500 106976 192506
rect 106924 192442 106976 192448
rect 107672 191282 107700 238726
rect 108592 231130 108620 239822
rect 109880 231198 109908 239822
rect 110616 238754 110644 240037
rect 111248 239850 111276 240037
rect 111892 239850 111920 240037
rect 110432 238726 110644 238754
rect 111168 239822 111276 239850
rect 111812 239822 111920 239850
rect 109868 231192 109920 231198
rect 109868 231134 109920 231140
rect 108580 231124 108632 231130
rect 108580 231066 108632 231072
rect 107660 191276 107712 191282
rect 107660 191218 107712 191224
rect 102140 191140 102192 191146
rect 102140 191082 102192 191088
rect 106188 189100 106240 189106
rect 106188 189042 106240 189048
rect 100668 186448 100720 186454
rect 100668 186390 100720 186396
rect 99286 183696 99342 183705
rect 99286 183631 99342 183640
rect 93860 182912 93912 182918
rect 93860 182854 93912 182860
rect 97540 182300 97592 182306
rect 97540 182242 97592 182248
rect 97552 177721 97580 182242
rect 99300 177721 99328 183631
rect 97538 177712 97594 177721
rect 97538 177647 97594 177656
rect 99286 177712 99342 177721
rect 99286 177647 99342 177656
rect 82820 177336 82872 177342
rect 82820 177278 82872 177284
rect 100680 176769 100708 186390
rect 106200 177721 106228 189042
rect 107568 187808 107620 187814
rect 107568 187750 107620 187756
rect 107580 177721 107608 187750
rect 110432 186998 110460 238726
rect 111168 219434 111196 239822
rect 111812 231198 111840 239822
rect 112548 235958 112576 240037
rect 113192 238754 113220 240037
rect 113192 238726 113404 238754
rect 113836 238746 113864 240037
rect 112536 235952 112588 235958
rect 112536 235894 112588 235900
rect 111800 231192 111852 231198
rect 111800 231134 111852 231140
rect 113376 220114 113404 238726
rect 113824 238740 113876 238746
rect 113824 238682 113876 238688
rect 114480 237318 114508 240037
rect 114560 239828 114612 239834
rect 114560 239770 114612 239776
rect 114468 237312 114520 237318
rect 114468 237254 114520 237260
rect 113364 220108 113416 220114
rect 113364 220050 113416 220056
rect 110524 219406 111196 219434
rect 110524 211886 110552 219406
rect 114572 213217 114600 239770
rect 115124 238542 115152 240037
rect 115756 239834 115784 240037
rect 115744 239828 115796 239834
rect 115744 239770 115796 239776
rect 116412 238754 116440 240037
rect 115952 238726 116440 238754
rect 115112 238536 115164 238542
rect 115112 238478 115164 238484
rect 114836 238196 114888 238202
rect 114836 238138 114888 238144
rect 114848 233238 114876 238138
rect 114836 233232 114888 233238
rect 114836 233174 114888 233180
rect 115952 220182 115980 238726
rect 117056 238678 117084 240037
rect 117044 238672 117096 238678
rect 117044 238614 117096 238620
rect 117700 235278 117728 240037
rect 118344 239970 118372 240037
rect 118332 239964 118384 239970
rect 118332 239906 118384 239912
rect 118988 239873 119016 240037
rect 118974 239864 119030 239873
rect 118974 239799 119030 239808
rect 119724 238754 119752 240094
rect 118712 238726 119752 238754
rect 117688 235272 117740 235278
rect 117688 235214 117740 235220
rect 115940 220176 115992 220182
rect 115940 220118 115992 220124
rect 114558 213208 114614 213217
rect 114558 213143 114614 213152
rect 110512 211880 110564 211886
rect 110512 211822 110564 211828
rect 110420 186992 110472 186998
rect 110420 186934 110472 186940
rect 118608 186380 118660 186386
rect 118608 186322 118660 186328
rect 114468 183592 114520 183598
rect 114468 183534 114520 183540
rect 112996 180872 113048 180878
rect 112996 180814 113048 180820
rect 110694 179480 110750 179489
rect 110694 179415 110750 179424
rect 109960 178084 110012 178090
rect 109960 178026 110012 178032
rect 106186 177712 106242 177721
rect 106186 177647 106242 177656
rect 107566 177712 107622 177721
rect 107566 177647 107622 177656
rect 104624 176996 104676 177002
rect 104624 176938 104676 176944
rect 103336 176928 103388 176934
rect 103336 176870 103388 176876
rect 103348 176769 103376 176870
rect 104636 176769 104664 176938
rect 109972 176769 110000 178026
rect 110708 177041 110736 179415
rect 113008 177177 113036 180814
rect 114480 177721 114508 183534
rect 116952 182368 117004 182374
rect 116952 182310 117004 182316
rect 115848 178152 115900 178158
rect 115848 178094 115900 178100
rect 114466 177712 114522 177721
rect 114466 177647 114522 177656
rect 112994 177168 113050 177177
rect 112994 177103 113050 177112
rect 110694 177032 110750 177041
rect 110694 176967 110750 176976
rect 115860 176769 115888 178094
rect 116964 177721 116992 182310
rect 118620 177721 118648 186322
rect 118712 185910 118740 238726
rect 119816 220250 119844 240887
rect 119804 220244 119856 220250
rect 119804 220186 119856 220192
rect 120092 202842 120120 250951
rect 120184 247625 120212 315250
rect 120276 261225 120304 324906
rect 121460 318776 121512 318782
rect 121460 318718 121512 318724
rect 121472 283778 121500 318718
rect 121552 309800 121604 309806
rect 121552 309742 121604 309748
rect 121564 291825 121592 309742
rect 122104 308440 122156 308446
rect 122104 308382 122156 308388
rect 121644 301504 121696 301510
rect 121644 301446 121696 301452
rect 121550 291816 121606 291825
rect 121550 291751 121606 291760
rect 121550 290456 121606 290465
rect 121550 290391 121606 290400
rect 121564 289950 121592 290391
rect 121552 289944 121604 289950
rect 121552 289886 121604 289892
rect 121552 289808 121604 289814
rect 121550 289776 121552 289785
rect 121604 289776 121606 289785
rect 121550 289711 121606 289720
rect 121550 288416 121606 288425
rect 121550 288351 121606 288360
rect 121564 287094 121592 288351
rect 121552 287088 121604 287094
rect 121552 287030 121604 287036
rect 121656 286385 121684 301446
rect 121734 291136 121790 291145
rect 121734 291071 121790 291080
rect 121748 289882 121776 291071
rect 121736 289876 121788 289882
rect 121736 289818 121788 289824
rect 122010 289096 122066 289105
rect 122010 289031 122066 289040
rect 121642 286376 121698 286385
rect 122024 286346 122052 289031
rect 122116 287065 122144 308382
rect 122102 287056 122158 287065
rect 122102 286991 122158 287000
rect 121642 286311 121698 286320
rect 122012 286340 122064 286346
rect 122012 286282 122064 286288
rect 122286 285696 122342 285705
rect 122286 285631 122342 285640
rect 121644 285592 121696 285598
rect 121644 285534 121696 285540
rect 121550 285016 121606 285025
rect 121550 284951 121606 284960
rect 121564 284374 121592 284951
rect 121552 284368 121604 284374
rect 121656 284345 121684 285534
rect 121552 284310 121604 284316
rect 121642 284336 121698 284345
rect 121642 284271 121698 284280
rect 121644 284232 121696 284238
rect 121644 284174 121696 284180
rect 121472 283750 121592 283778
rect 121458 282976 121514 282985
rect 121458 282911 121460 282920
rect 121512 282911 121514 282920
rect 121460 282882 121512 282888
rect 121460 281648 121512 281654
rect 121458 281616 121460 281625
rect 121512 281616 121514 281625
rect 121458 281551 121514 281560
rect 121460 280288 121512 280294
rect 121458 280256 121460 280265
rect 121512 280256 121514 280265
rect 121458 280191 121514 280200
rect 121458 278896 121514 278905
rect 121458 278831 121460 278840
rect 121512 278831 121514 278840
rect 121460 278802 121512 278808
rect 121458 277536 121514 277545
rect 121458 277471 121514 277480
rect 121472 277438 121500 277471
rect 121460 277432 121512 277438
rect 121460 277374 121512 277380
rect 121458 276856 121514 276865
rect 121458 276791 121514 276800
rect 121472 276078 121500 276791
rect 121460 276072 121512 276078
rect 121460 276014 121512 276020
rect 121458 274816 121514 274825
rect 121458 274751 121514 274760
rect 121472 274718 121500 274751
rect 121460 274712 121512 274718
rect 121460 274654 121512 274660
rect 121460 274304 121512 274310
rect 121460 274246 121512 274252
rect 121472 274145 121500 274246
rect 121458 274136 121514 274145
rect 121458 274071 121514 274080
rect 121458 273456 121514 273465
rect 121458 273391 121514 273400
rect 121472 273290 121500 273391
rect 121460 273284 121512 273290
rect 121460 273226 121512 273232
rect 121564 272785 121592 283750
rect 121656 283665 121684 284174
rect 121642 283656 121698 283665
rect 121642 283591 121698 283600
rect 121642 282296 121698 282305
rect 121642 282231 121698 282240
rect 121656 281586 121684 282231
rect 121644 281580 121696 281586
rect 121644 281522 121696 281528
rect 121642 280936 121698 280945
rect 121642 280871 121698 280880
rect 121656 280226 121684 280871
rect 121644 280220 121696 280226
rect 121644 280162 121696 280168
rect 121642 279576 121698 279585
rect 121642 279511 121698 279520
rect 121656 278798 121684 279511
rect 121644 278792 121696 278798
rect 121644 278734 121696 278740
rect 121642 278216 121698 278225
rect 121642 278151 121698 278160
rect 121656 277506 121684 278151
rect 121644 277500 121696 277506
rect 121644 277442 121696 277448
rect 121642 276176 121698 276185
rect 121642 276111 121698 276120
rect 121550 272776 121606 272785
rect 121550 272711 121606 272720
rect 121550 271416 121606 271425
rect 121550 271351 121606 271360
rect 121458 270056 121514 270065
rect 121458 269991 121514 270000
rect 121472 269142 121500 269991
rect 121460 269136 121512 269142
rect 121460 269078 121512 269084
rect 121564 268394 121592 271351
rect 121656 271182 121684 276111
rect 122102 275496 122158 275505
rect 122102 275431 122158 275440
rect 121644 271176 121696 271182
rect 121644 271118 121696 271124
rect 121552 268388 121604 268394
rect 121552 268330 121604 268336
rect 121458 268016 121514 268025
rect 121458 267951 121514 267960
rect 121472 267782 121500 267951
rect 121460 267776 121512 267782
rect 121460 267718 121512 267724
rect 121550 267336 121606 267345
rect 121550 267271 121606 267280
rect 121458 266656 121514 266665
rect 121458 266591 121514 266600
rect 121472 266490 121500 266591
rect 121460 266484 121512 266490
rect 121460 266426 121512 266432
rect 121564 266422 121592 267271
rect 121644 267028 121696 267034
rect 121644 266970 121696 266976
rect 121552 266416 121604 266422
rect 121552 266358 121604 266364
rect 121550 265976 121606 265985
rect 121550 265911 121606 265920
rect 121458 265296 121514 265305
rect 121458 265231 121514 265240
rect 121472 265062 121500 265231
rect 121460 265056 121512 265062
rect 121460 264998 121512 265004
rect 121564 264994 121592 265911
rect 121552 264988 121604 264994
rect 121552 264930 121604 264936
rect 121656 264625 121684 266970
rect 121642 264616 121698 264625
rect 121642 264551 121698 264560
rect 122116 264217 122144 275431
rect 122300 275330 122328 285631
rect 122288 275324 122340 275330
rect 122288 275266 122340 275272
rect 122102 264208 122158 264217
rect 122102 264143 122158 264152
rect 121550 263936 121606 263945
rect 121550 263871 121606 263880
rect 121564 263634 121592 263871
rect 121552 263628 121604 263634
rect 121552 263570 121604 263576
rect 121460 263560 121512 263566
rect 121460 263502 121512 263508
rect 121472 263265 121500 263502
rect 121458 263256 121514 263265
rect 121458 263191 121514 263200
rect 121458 262576 121514 262585
rect 121458 262511 121514 262520
rect 121472 262274 121500 262511
rect 121460 262268 121512 262274
rect 121460 262210 121512 262216
rect 121458 261896 121514 261905
rect 121458 261831 121514 261840
rect 120262 261216 120318 261225
rect 120262 261151 120318 261160
rect 121472 260914 121500 261831
rect 121460 260908 121512 260914
rect 121460 260850 121512 260856
rect 121458 259856 121514 259865
rect 121458 259791 121514 259800
rect 121472 259486 121500 259791
rect 121460 259480 121512 259486
rect 121460 259422 121512 259428
rect 121552 259412 121604 259418
rect 121552 259354 121604 259360
rect 121458 259176 121514 259185
rect 121458 259111 121514 259120
rect 121472 258126 121500 259111
rect 121564 258505 121592 259354
rect 121550 258496 121606 258505
rect 121550 258431 121606 258440
rect 121460 258120 121512 258126
rect 121460 258062 121512 258068
rect 121460 257916 121512 257922
rect 121460 257858 121512 257864
rect 121472 257145 121500 257858
rect 121550 257816 121606 257825
rect 121550 257751 121606 257760
rect 121458 257136 121514 257145
rect 121458 257071 121514 257080
rect 121564 256766 121592 257751
rect 121552 256760 121604 256766
rect 121552 256702 121604 256708
rect 121644 256692 121696 256698
rect 121644 256634 121696 256640
rect 121460 256624 121512 256630
rect 121460 256566 121512 256572
rect 121472 256465 121500 256566
rect 121458 256456 121514 256465
rect 121458 256391 121514 256400
rect 121656 255785 121684 256634
rect 121642 255776 121698 255785
rect 121642 255711 121698 255720
rect 121550 255096 121606 255105
rect 121550 255031 121606 255040
rect 121458 254416 121514 254425
rect 121458 254351 121514 254360
rect 121472 254046 121500 254351
rect 121460 254040 121512 254046
rect 121460 253982 121512 253988
rect 121564 253978 121592 255031
rect 121552 253972 121604 253978
rect 121552 253914 121604 253920
rect 122102 253736 122158 253745
rect 122102 253671 122158 253680
rect 121550 253056 121606 253065
rect 121550 252991 121606 253000
rect 121564 252618 121592 252991
rect 121552 252612 121604 252618
rect 121552 252554 121604 252560
rect 121460 252544 121512 252550
rect 121460 252486 121512 252492
rect 121472 252385 121500 252486
rect 121458 252376 121514 252385
rect 121458 252311 121514 252320
rect 121458 251696 121514 251705
rect 121458 251631 121514 251640
rect 121472 250510 121500 251631
rect 121460 250504 121512 250510
rect 121460 250446 121512 250452
rect 121550 250336 121606 250345
rect 121550 250271 121606 250280
rect 121564 249830 121592 250271
rect 121552 249824 121604 249830
rect 121552 249766 121604 249772
rect 121460 249756 121512 249762
rect 121460 249698 121512 249704
rect 121472 249665 121500 249698
rect 121458 249656 121514 249665
rect 121458 249591 121514 249600
rect 121458 248976 121514 248985
rect 121458 248911 121514 248920
rect 121472 248470 121500 248911
rect 121460 248464 121512 248470
rect 121460 248406 121512 248412
rect 121458 248296 121514 248305
rect 121458 248231 121514 248240
rect 120170 247616 120226 247625
rect 120170 247551 120226 247560
rect 121472 247110 121500 248231
rect 121460 247104 121512 247110
rect 121460 247046 121512 247052
rect 121550 246936 121606 246945
rect 121550 246871 121606 246880
rect 121564 245682 121592 246871
rect 121552 245676 121604 245682
rect 121552 245618 121604 245624
rect 121460 245608 121512 245614
rect 121460 245550 121512 245556
rect 121550 245576 121606 245585
rect 121472 244905 121500 245550
rect 121550 245511 121606 245520
rect 121458 244896 121514 244905
rect 121458 244831 121514 244840
rect 121564 244390 121592 245511
rect 121552 244384 121604 244390
rect 121552 244326 121604 244332
rect 121460 244248 121512 244254
rect 121460 244190 121512 244196
rect 121642 244216 121698 244225
rect 121472 243545 121500 244190
rect 121642 244151 121698 244160
rect 121458 243536 121514 243545
rect 121458 243471 121514 243480
rect 121552 242888 121604 242894
rect 121458 242856 121514 242865
rect 121552 242830 121604 242836
rect 121458 242791 121460 242800
rect 121512 242791 121514 242800
rect 121460 242762 121512 242768
rect 121564 242185 121592 242830
rect 121656 242214 121684 244151
rect 122116 243574 122144 253671
rect 122104 243568 122156 243574
rect 122104 243510 122156 243516
rect 121644 242208 121696 242214
rect 121550 242176 121606 242185
rect 121644 242150 121696 242156
rect 121550 242111 121606 242120
rect 121458 240816 121514 240825
rect 121458 240751 121514 240760
rect 121472 240242 121500 240751
rect 121460 240236 121512 240242
rect 121460 240178 121512 240184
rect 121552 240168 121604 240174
rect 121550 240136 121552 240145
rect 121604 240136 121606 240145
rect 121550 240071 121606 240080
rect 123496 239970 123524 643078
rect 123576 536852 123628 536858
rect 123576 536794 123628 536800
rect 123484 239964 123536 239970
rect 123484 239906 123536 239912
rect 123588 238542 123616 536794
rect 123668 309800 123720 309806
rect 123668 309742 123720 309748
rect 123680 274310 123708 309742
rect 124876 284238 124904 702578
rect 126244 683188 126296 683194
rect 126244 683130 126296 683136
rect 124956 470620 125008 470626
rect 124956 470562 125008 470568
rect 124968 285598 124996 470562
rect 125048 312588 125100 312594
rect 125048 312530 125100 312536
rect 124956 285592 125008 285598
rect 124956 285534 125008 285540
rect 124864 284232 124916 284238
rect 124864 284174 124916 284180
rect 123668 274304 123720 274310
rect 123668 274246 123720 274252
rect 125060 257922 125088 312530
rect 125600 293276 125652 293282
rect 125600 293218 125652 293224
rect 125612 263566 125640 293218
rect 125600 263560 125652 263566
rect 125600 263502 125652 263508
rect 125048 257916 125100 257922
rect 125048 257858 125100 257864
rect 124864 257372 124916 257378
rect 124864 257314 124916 257320
rect 124876 238678 124904 257314
rect 126256 252550 126284 683130
rect 126336 484424 126388 484430
rect 126336 484366 126388 484372
rect 126348 267034 126376 484366
rect 127624 378208 127676 378214
rect 127624 378150 127676 378156
rect 127636 289814 127664 378150
rect 127714 292768 127770 292777
rect 127714 292703 127770 292712
rect 127624 289808 127676 289814
rect 127624 289750 127676 289756
rect 126336 267028 126388 267034
rect 126336 266970 126388 266976
rect 126244 252544 126296 252550
rect 126244 252486 126296 252492
rect 124864 238672 124916 238678
rect 124864 238614 124916 238620
rect 123576 238536 123628 238542
rect 123576 238478 123628 238484
rect 127728 206990 127756 292703
rect 129016 245614 129044 702850
rect 133144 702568 133196 702574
rect 133144 702510 133196 702516
rect 130384 616888 130436 616894
rect 130384 616830 130436 616836
rect 129096 430636 129148 430642
rect 129096 430578 129148 430584
rect 129108 256630 129136 430578
rect 130396 256698 130424 616830
rect 130476 271924 130528 271930
rect 130476 271866 130528 271872
rect 130384 256692 130436 256698
rect 130384 256634 130436 256640
rect 129096 256624 129148 256630
rect 129096 256566 129148 256572
rect 129004 245608 129056 245614
rect 129004 245550 129056 245556
rect 128360 244316 128412 244322
rect 128360 244258 128412 244264
rect 128372 242826 128400 244258
rect 128360 242820 128412 242826
rect 128360 242762 128412 242768
rect 130488 238610 130516 271866
rect 133156 242894 133184 702510
rect 137848 697678 137876 703520
rect 154132 700330 154160 703520
rect 170324 702434 170352 703520
rect 202800 703118 202828 703520
rect 201500 703112 201552 703118
rect 201500 703054 201552 703060
rect 202788 703112 202840 703118
rect 202788 703054 202840 703060
rect 169772 702406 170352 702434
rect 154120 700324 154172 700330
rect 154120 700266 154172 700272
rect 151084 698964 151136 698970
rect 151084 698906 151136 698912
rect 137836 697672 137888 697678
rect 137836 697614 137888 697620
rect 134524 697604 134576 697610
rect 134524 697546 134576 697552
rect 134536 244254 134564 697546
rect 148324 670744 148376 670750
rect 148324 670686 148376 670692
rect 142804 576904 142856 576910
rect 142804 576846 142856 576852
rect 141424 524476 141476 524482
rect 141424 524418 141476 524424
rect 137284 294228 137336 294234
rect 137284 294170 137336 294176
rect 134524 244248 134576 244254
rect 134524 244190 134576 244196
rect 133144 242888 133196 242894
rect 133144 242830 133196 242836
rect 130476 238604 130528 238610
rect 130476 238546 130528 238552
rect 137296 217462 137324 294170
rect 141436 249762 141464 524418
rect 142816 253201 142844 576846
rect 148336 319462 148364 670686
rect 148324 319456 148376 319462
rect 148324 319398 148376 319404
rect 148324 298512 148376 298518
rect 148324 298454 148376 298460
rect 146944 295724 146996 295730
rect 146944 295666 146996 295672
rect 144184 276072 144236 276078
rect 144184 276014 144236 276020
rect 144196 262886 144224 276014
rect 144184 262880 144236 262886
rect 144184 262822 144236 262828
rect 142802 253192 142858 253201
rect 142802 253127 142858 253136
rect 141424 249756 141476 249762
rect 141424 249698 141476 249704
rect 137284 217456 137336 217462
rect 137284 217398 137336 217404
rect 146956 210526 146984 295666
rect 146944 210520 146996 210526
rect 146944 210462 146996 210468
rect 127716 206984 127768 206990
rect 127716 206926 127768 206932
rect 148336 205018 148364 298454
rect 151096 259418 151124 698906
rect 169772 305658 169800 702406
rect 201512 308446 201540 703054
rect 218992 699718 219020 703520
rect 214564 699712 214616 699718
rect 214564 699654 214616 699660
rect 218980 699712 219032 699718
rect 218980 699654 219032 699660
rect 201500 308440 201552 308446
rect 201500 308382 201552 308388
rect 169760 305652 169812 305658
rect 169760 305594 169812 305600
rect 170404 303816 170456 303822
rect 170404 303758 170456 303764
rect 169024 297084 169076 297090
rect 169024 297026 169076 297032
rect 152464 294296 152516 294302
rect 152464 294238 152516 294244
rect 151084 259412 151136 259418
rect 151084 259354 151136 259360
rect 148324 205012 148376 205018
rect 148324 204954 148376 204960
rect 120080 202836 120132 202842
rect 120080 202778 120132 202784
rect 133788 187740 133840 187746
rect 133788 187682 133840 187688
rect 132408 186516 132460 186522
rect 132408 186458 132460 186464
rect 118700 185904 118752 185910
rect 118700 185846 118752 185852
rect 121368 184952 121420 184958
rect 121368 184894 121420 184900
rect 121380 177721 121408 184894
rect 129464 182232 129516 182238
rect 129464 182174 129516 182180
rect 123760 179512 123812 179518
rect 123760 179454 123812 179460
rect 116950 177712 117006 177721
rect 116950 177647 117006 177656
rect 118606 177712 118662 177721
rect 118606 177647 118662 177656
rect 121366 177712 121422 177721
rect 121366 177647 121422 177656
rect 123772 177041 123800 179454
rect 128084 179444 128136 179450
rect 128084 179386 128136 179392
rect 126060 178220 126112 178226
rect 126060 178162 126112 178168
rect 123758 177032 123814 177041
rect 123758 176967 123814 176976
rect 124496 176792 124548 176798
rect 100666 176760 100722 176769
rect 100666 176695 100722 176704
rect 103334 176760 103390 176769
rect 103334 176695 103390 176704
rect 104622 176760 104678 176769
rect 104622 176695 104678 176704
rect 108118 176760 108174 176769
rect 108118 176695 108120 176704
rect 108172 176695 108174 176704
rect 109958 176760 110014 176769
rect 109958 176695 110014 176704
rect 115846 176760 115902 176769
rect 115846 176695 115902 176704
rect 124494 176760 124496 176769
rect 126072 176769 126100 178162
rect 128096 177041 128124 179386
rect 129476 177721 129504 182174
rect 132420 177721 132448 186458
rect 133800 177721 133828 187682
rect 152476 186998 152504 294238
rect 162124 292868 162176 292874
rect 162124 292810 162176 292816
rect 160744 292800 160796 292806
rect 160744 292742 160796 292748
rect 155224 291372 155276 291378
rect 155224 291314 155276 291320
rect 155236 203590 155264 291314
rect 160756 242282 160784 292742
rect 160744 242276 160796 242282
rect 160744 242218 160796 242224
rect 160744 231260 160796 231266
rect 160744 231202 160796 231208
rect 155224 203584 155276 203590
rect 155224 203526 155276 203532
rect 160756 188630 160784 231202
rect 160744 188624 160796 188630
rect 160744 188566 160796 188572
rect 152464 186992 152516 186998
rect 152464 186934 152516 186940
rect 162136 178702 162164 292810
rect 169036 189854 169064 297026
rect 169024 189848 169076 189854
rect 169024 189790 169076 189796
rect 169024 186448 169076 186454
rect 169024 186390 169076 186396
rect 167736 182368 167788 182374
rect 167736 182310 167788 182316
rect 166356 180872 166408 180878
rect 166356 180814 166408 180820
rect 162124 178696 162176 178702
rect 162124 178638 162176 178644
rect 148232 178356 148284 178362
rect 148232 178298 148284 178304
rect 134800 178288 134852 178294
rect 134800 178230 134852 178236
rect 129462 177712 129518 177721
rect 129462 177647 129518 177656
rect 132406 177712 132462 177721
rect 132406 177647 132462 177656
rect 133786 177712 133842 177721
rect 133786 177647 133842 177656
rect 130752 177064 130804 177070
rect 128082 177032 128138 177041
rect 130752 177006 130804 177012
rect 128082 176967 128138 176976
rect 130764 176769 130792 177006
rect 134812 176769 134840 178230
rect 136088 176860 136140 176866
rect 136088 176802 136140 176808
rect 136100 176769 136128 176802
rect 148244 176769 148272 178298
rect 165344 178288 165396 178294
rect 165344 178230 165396 178236
rect 124548 176760 124550 176769
rect 124494 176695 124550 176704
rect 126058 176760 126114 176769
rect 126058 176695 126114 176704
rect 130750 176760 130806 176769
rect 130750 176695 130806 176704
rect 134798 176760 134854 176769
rect 134798 176695 134854 176704
rect 136086 176760 136142 176769
rect 136086 176695 136142 176704
rect 148230 176760 148286 176769
rect 148230 176695 148286 176704
rect 108120 176666 108172 176672
rect 158904 176316 158956 176322
rect 158904 176258 158956 176264
rect 121920 176248 121972 176254
rect 121920 176190 121972 176196
rect 113180 176180 113232 176186
rect 113180 176122 113232 176128
rect 100760 175976 100812 175982
rect 100760 175918 100812 175924
rect 100772 175409 100800 175918
rect 100758 175400 100814 175409
rect 100758 175335 100814 175344
rect 113192 175001 113220 176122
rect 119436 176044 119488 176050
rect 119436 175986 119488 175992
rect 119448 175001 119476 175986
rect 121932 175409 121960 176190
rect 128176 176112 128228 176118
rect 128176 176054 128228 176060
rect 128188 175409 128216 176054
rect 158916 175409 158944 176258
rect 121918 175400 121974 175409
rect 121918 175335 121974 175344
rect 128174 175400 128230 175409
rect 128174 175335 128230 175344
rect 158902 175400 158958 175409
rect 158902 175335 158958 175344
rect 165356 175234 165384 178230
rect 165528 177064 165580 177070
rect 165528 177006 165580 177012
rect 165436 176996 165488 177002
rect 165436 176938 165488 176944
rect 165344 175228 165396 175234
rect 165344 175170 165396 175176
rect 113178 174992 113234 175001
rect 113178 174927 113234 174936
rect 119434 174992 119490 175001
rect 119434 174927 119490 174936
rect 165448 173194 165476 176938
rect 165540 174554 165568 177006
rect 166264 176316 166316 176322
rect 166264 176258 166316 176264
rect 165528 174548 165580 174554
rect 165528 174490 165580 174496
rect 165436 173188 165488 173194
rect 165436 173130 165488 173136
rect 166276 149054 166304 176258
rect 166368 164218 166396 180814
rect 166448 178152 166500 178158
rect 166448 178094 166500 178100
rect 166460 165578 166488 178094
rect 167644 176928 167696 176934
rect 167644 176870 167696 176876
rect 166540 176248 166592 176254
rect 166540 176190 166592 176196
rect 166552 168366 166580 176190
rect 166540 168360 166592 168366
rect 166540 168302 166592 168308
rect 166448 165572 166500 165578
rect 166448 165514 166500 165520
rect 166356 164212 166408 164218
rect 166356 164154 166408 164160
rect 167656 158710 167684 176870
rect 167748 167006 167776 182310
rect 167828 179512 167880 179518
rect 167828 179454 167880 179460
rect 167840 169726 167868 179454
rect 167920 178220 167972 178226
rect 167920 178162 167972 178168
rect 167932 171086 167960 178162
rect 168010 171592 168066 171601
rect 168010 171527 168066 171536
rect 168024 171154 168052 171527
rect 168012 171148 168064 171154
rect 168012 171090 168064 171096
rect 167920 171080 167972 171086
rect 167920 171022 167972 171028
rect 167828 169720 167880 169726
rect 167828 169662 167880 169668
rect 167736 167000 167788 167006
rect 167736 166942 167788 166948
rect 167644 158704 167696 158710
rect 167644 158646 167696 158652
rect 169036 157350 169064 186390
rect 169300 183592 169352 183598
rect 169300 183534 169352 183540
rect 169208 182300 169260 182306
rect 169208 182242 169260 182248
rect 169116 178356 169168 178362
rect 169116 178298 169168 178304
rect 169024 157344 169076 157350
rect 169024 157286 169076 157292
rect 169128 150414 169156 178298
rect 169220 155922 169248 182242
rect 169312 165510 169340 183534
rect 170416 181558 170444 303758
rect 213184 302456 213236 302462
rect 213184 302398 213236 302404
rect 206284 299736 206336 299742
rect 206284 299678 206336 299684
rect 202144 299668 202196 299674
rect 202144 299610 202196 299616
rect 186964 298444 187016 298450
rect 186964 298386 187016 298392
rect 177302 294264 177358 294273
rect 177302 294199 177358 294208
rect 173164 189100 173216 189106
rect 173164 189042 173216 189048
rect 171784 187808 171836 187814
rect 171784 187750 171836 187756
rect 170588 186516 170640 186522
rect 170588 186458 170640 186464
rect 170496 184952 170548 184958
rect 170496 184894 170548 184900
rect 170404 181552 170456 181558
rect 170404 181494 170456 181500
rect 170404 178084 170456 178090
rect 170404 178026 170456 178032
rect 169300 165504 169352 165510
rect 169300 165446 169352 165452
rect 170416 162858 170444 178026
rect 170508 168298 170536 184894
rect 170600 173874 170628 186458
rect 170680 176180 170732 176186
rect 170680 176122 170732 176128
rect 170588 173868 170640 173874
rect 170588 173810 170640 173816
rect 170496 168292 170548 168298
rect 170496 168234 170548 168240
rect 170692 164150 170720 176122
rect 170680 164144 170732 164150
rect 170680 164086 170732 164092
rect 170404 162852 170456 162858
rect 170404 162794 170456 162800
rect 171796 161430 171824 187750
rect 171784 161424 171836 161430
rect 171784 161366 171836 161372
rect 173176 160070 173204 189042
rect 173164 160064 173216 160070
rect 173164 160006 173216 160012
rect 169208 155916 169260 155922
rect 169208 155858 169260 155864
rect 173256 151088 173308 151094
rect 173256 151030 173308 151036
rect 169116 150408 169168 150414
rect 169116 150350 169168 150356
rect 166264 149048 166316 149054
rect 166264 148990 166316 148996
rect 167736 147688 167788 147694
rect 167736 147630 167788 147636
rect 166264 143608 166316 143614
rect 166264 143550 166316 143556
rect 66166 129296 66222 129305
rect 66166 129231 66222 129240
rect 65154 126304 65210 126313
rect 65154 126239 65210 126248
rect 65168 125662 65196 126239
rect 62028 125656 62080 125662
rect 62028 125598 62080 125604
rect 65156 125656 65208 125662
rect 65156 125598 65208 125604
rect 62040 93838 62068 125598
rect 66074 125216 66130 125225
rect 66074 125151 66130 125160
rect 65982 123584 66038 123593
rect 65982 123519 66038 123528
rect 65996 122913 66024 123519
rect 64786 122904 64842 122913
rect 64786 122839 64842 122848
rect 65982 122904 66038 122913
rect 65982 122839 66038 122848
rect 62028 93832 62080 93838
rect 62028 93774 62080 93780
rect 64800 89690 64828 122839
rect 65982 122632 66038 122641
rect 65982 122567 66038 122576
rect 65996 91089 66024 122567
rect 65982 91080 66038 91089
rect 66088 91050 66116 125151
rect 66180 94897 66208 129231
rect 67546 128072 67602 128081
rect 67546 128007 67602 128016
rect 67454 120864 67510 120873
rect 67454 120799 67510 120808
rect 67362 102368 67418 102377
rect 67362 102303 67418 102312
rect 66166 94888 66222 94897
rect 66166 94823 66222 94832
rect 65982 91015 66038 91024
rect 66076 91044 66128 91050
rect 66076 90986 66128 90992
rect 64788 89684 64840 89690
rect 64788 89626 64840 89632
rect 67376 85542 67404 102303
rect 67468 88262 67496 120799
rect 67560 93809 67588 128007
rect 67638 100736 67694 100745
rect 67638 100671 67694 100680
rect 67546 93800 67602 93809
rect 67546 93735 67602 93744
rect 67652 88330 67680 100671
rect 164976 98048 165028 98054
rect 164976 97990 165028 97996
rect 164882 95160 164938 95169
rect 164882 95095 164938 95104
rect 111982 94752 112038 94761
rect 111982 94687 112038 94696
rect 113730 94752 113786 94761
rect 113730 94687 113786 94696
rect 129370 94752 129426 94761
rect 129370 94687 129426 94696
rect 151634 94752 151690 94761
rect 151634 94687 151690 94696
rect 111996 93974 112024 94687
rect 111984 93968 112036 93974
rect 111984 93910 112036 93916
rect 113744 93906 113772 94687
rect 122840 94512 122892 94518
rect 122840 94454 122892 94460
rect 113732 93900 113784 93906
rect 113732 93842 113784 93848
rect 118054 93664 118110 93673
rect 118054 93599 118110 93608
rect 85670 93528 85726 93537
rect 85670 93463 85726 93472
rect 107750 93528 107806 93537
rect 107750 93463 107806 93472
rect 85684 93158 85712 93463
rect 107764 93226 107792 93463
rect 118068 93362 118096 93599
rect 120630 93528 120686 93537
rect 120630 93463 120686 93472
rect 118056 93356 118108 93362
rect 118056 93298 118108 93304
rect 120644 93294 120672 93463
rect 120632 93288 120684 93294
rect 110142 93256 110198 93265
rect 107752 93220 107804 93226
rect 120632 93230 120684 93236
rect 110142 93191 110198 93200
rect 107752 93162 107804 93168
rect 85672 93152 85724 93158
rect 85672 93094 85724 93100
rect 85118 92440 85174 92449
rect 85118 92375 85174 92384
rect 91650 92440 91706 92449
rect 91650 92375 91706 92384
rect 95054 92440 95110 92449
rect 95054 92375 95056 92384
rect 75826 91216 75882 91225
rect 75826 91151 75882 91160
rect 67640 88324 67692 88330
rect 67640 88266 67692 88272
rect 67456 88256 67508 88262
rect 67456 88198 67508 88204
rect 67364 85536 67416 85542
rect 67364 85478 67416 85484
rect 75840 77246 75868 91151
rect 85132 91118 85160 92375
rect 90638 91760 90694 91769
rect 90638 91695 90694 91704
rect 86866 91216 86922 91225
rect 86866 91151 86922 91160
rect 88062 91216 88118 91225
rect 88062 91151 88118 91160
rect 89626 91216 89682 91225
rect 89626 91151 89682 91160
rect 85120 91112 85172 91118
rect 85120 91054 85172 91060
rect 86880 84046 86908 91151
rect 88076 86902 88104 91151
rect 88064 86896 88116 86902
rect 88064 86838 88116 86844
rect 86868 84040 86920 84046
rect 86868 83982 86920 83988
rect 89640 82754 89668 91151
rect 90652 89622 90680 91695
rect 91664 91186 91692 92375
rect 95108 92375 95110 92384
rect 106002 92440 106058 92449
rect 106002 92375 106058 92384
rect 95056 92346 95108 92352
rect 102690 91760 102746 91769
rect 102690 91695 102746 91704
rect 100022 91624 100078 91633
rect 100022 91559 100078 91568
rect 99286 91488 99342 91497
rect 99286 91423 99342 91432
rect 97814 91352 97870 91361
rect 97814 91287 97870 91296
rect 99102 91352 99158 91361
rect 99102 91287 99158 91296
rect 93766 91216 93822 91225
rect 91652 91180 91704 91186
rect 93766 91151 93822 91160
rect 95146 91216 95202 91225
rect 95146 91151 95202 91160
rect 96526 91216 96582 91225
rect 96526 91151 96582 91160
rect 91652 91122 91704 91128
rect 90640 89616 90692 89622
rect 90640 89558 90692 89564
rect 89628 82748 89680 82754
rect 89628 82690 89680 82696
rect 93780 81326 93808 91151
rect 93768 81320 93820 81326
rect 93768 81262 93820 81268
rect 95160 79898 95188 91151
rect 96540 83978 96568 91151
rect 96528 83972 96580 83978
rect 96528 83914 96580 83920
rect 97828 81433 97856 91287
rect 97906 91216 97962 91225
rect 97906 91151 97962 91160
rect 97814 81424 97870 81433
rect 97814 81359 97870 81368
rect 95148 79892 95200 79898
rect 95148 79834 95200 79840
rect 97920 78674 97948 91151
rect 99116 82686 99144 91287
rect 99194 91216 99250 91225
rect 99194 91151 99250 91160
rect 99104 82680 99156 82686
rect 99104 82622 99156 82628
rect 99208 80073 99236 91151
rect 99194 80064 99250 80073
rect 99194 79999 99250 80008
rect 97908 78668 97960 78674
rect 97908 78610 97960 78616
rect 99300 78577 99328 91423
rect 100036 89486 100064 91559
rect 101862 91488 101918 91497
rect 101862 91423 101918 91432
rect 100574 91216 100630 91225
rect 100574 91151 100630 91160
rect 100024 89480 100076 89486
rect 100024 89422 100076 89428
rect 100588 85338 100616 91151
rect 101876 86970 101904 91423
rect 102046 91352 102102 91361
rect 102046 91287 102102 91296
rect 101954 91216 102010 91225
rect 101954 91151 102010 91160
rect 101864 86964 101916 86970
rect 101864 86906 101916 86912
rect 100576 85332 100628 85338
rect 100576 85274 100628 85280
rect 101968 82550 101996 91151
rect 101956 82544 102008 82550
rect 101956 82486 102008 82492
rect 99286 78568 99342 78577
rect 102060 78538 102088 91287
rect 102704 89554 102732 91695
rect 104254 91216 104310 91225
rect 104254 91151 104310 91160
rect 104806 91216 104862 91225
rect 104806 91151 104862 91160
rect 102692 89548 102744 89554
rect 102692 89490 102744 89496
rect 104268 85406 104296 91151
rect 104256 85400 104308 85406
rect 104256 85342 104308 85348
rect 104820 84182 104848 91151
rect 106016 90914 106044 92375
rect 107566 91352 107622 91361
rect 107566 91287 107622 91296
rect 106186 91216 106242 91225
rect 106186 91151 106242 91160
rect 107474 91216 107530 91225
rect 107474 91151 107530 91160
rect 106004 90908 106056 90914
rect 106004 90850 106056 90856
rect 104808 84176 104860 84182
rect 104808 84118 104860 84124
rect 106200 83910 106228 91151
rect 106188 83904 106240 83910
rect 106188 83846 106240 83852
rect 107488 81190 107516 91151
rect 107476 81184 107528 81190
rect 107476 81126 107528 81132
rect 99286 78503 99342 78512
rect 102048 78532 102100 78538
rect 102048 78474 102100 78480
rect 75828 77240 75880 77246
rect 75828 77182 75880 77188
rect 82820 76560 82872 76566
rect 82820 76502 82872 76508
rect 56600 73840 56652 73846
rect 56600 73782 56652 73788
rect 53104 71732 53156 71738
rect 53104 71674 53156 71680
rect 52460 71052 52512 71058
rect 52460 70994 52512 71000
rect 51724 13184 51776 13190
rect 51724 13126 51776 13132
rect 51080 13116 51132 13122
rect 51080 13058 51132 13064
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51092 354 51120 13058
rect 52472 3534 52500 70994
rect 52552 35216 52604 35222
rect 52552 35158 52604 35164
rect 52460 3528 52512 3534
rect 52460 3470 52512 3476
rect 52564 480 52592 35158
rect 56612 16574 56640 73782
rect 64880 72480 64932 72486
rect 64880 72422 64932 72428
rect 60740 49020 60792 49026
rect 60740 48962 60792 48968
rect 57980 39432 58032 39438
rect 57980 39374 58032 39380
rect 57992 16574 58020 39374
rect 59358 30968 59414 30977
rect 59358 30903 59414 30912
rect 56612 16546 56824 16574
rect 57992 16546 58480 16574
rect 54942 13016 54998 13025
rect 54942 12951 54998 12960
rect 53380 3528 53432 3534
rect 53380 3470 53432 3476
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53392 354 53420 3470
rect 54956 480 54984 12951
rect 56048 4820 56100 4826
rect 56048 4762 56100 4768
rect 56060 480 56088 4762
rect 53718 354 53830 480
rect 53392 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58452 480 58480 16546
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 30903
rect 60752 16574 60780 48962
rect 63500 22772 63552 22778
rect 63500 22714 63552 22720
rect 63512 16574 63540 22714
rect 64892 16574 64920 72422
rect 69020 64252 69072 64258
rect 69020 64194 69072 64200
rect 66260 39364 66312 39370
rect 66260 39306 66312 39312
rect 66272 16574 66300 39306
rect 60752 16546 60872 16574
rect 63512 16546 64368 16574
rect 64892 16546 65104 16574
rect 66272 16546 66760 16574
rect 60844 480 60872 16546
rect 61568 14544 61620 14550
rect 61568 14486 61620 14492
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61580 354 61608 14486
rect 63224 3460 63276 3466
rect 63224 3402 63276 3408
rect 63236 480 63264 3402
rect 64340 480 64368 16546
rect 61998 354 62110 480
rect 61580 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66732 480 66760 16546
rect 67916 3596 67968 3602
rect 67916 3538 67968 3544
rect 67928 480 67956 3538
rect 69032 3534 69060 64194
rect 71780 62824 71832 62830
rect 71780 62766 71832 62772
rect 70400 58744 70452 58750
rect 70400 58686 70452 58692
rect 70412 16574 70440 58686
rect 71792 16574 71820 62766
rect 73160 55888 73212 55894
rect 73160 55830 73212 55836
rect 73172 16574 73200 55830
rect 81440 50380 81492 50386
rect 81440 50322 81492 50328
rect 80060 42152 80112 42158
rect 80060 42094 80112 42100
rect 77300 40792 77352 40798
rect 77300 40734 77352 40740
rect 75920 28348 75972 28354
rect 75920 28290 75972 28296
rect 70412 16546 71544 16574
rect 71792 16546 72648 16574
rect 73172 16546 73384 16574
rect 69112 15972 69164 15978
rect 69112 15914 69164 15920
rect 69020 3528 69072 3534
rect 69020 3470 69072 3476
rect 69124 480 69152 15914
rect 69940 3528 69992 3534
rect 69940 3470 69992 3476
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 69952 354 69980 3470
rect 71516 480 71544 16546
rect 72620 480 72648 16546
rect 70278 354 70390 480
rect 69952 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75000 8968 75052 8974
rect 75000 8910 75052 8916
rect 75012 480 75040 8910
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 28290
rect 77312 6914 77340 40734
rect 77390 29608 77446 29617
rect 77390 29543 77446 29552
rect 77404 16574 77432 29543
rect 78680 17332 78732 17338
rect 78680 17274 78732 17280
rect 78692 16574 78720 17274
rect 80072 16574 80100 42094
rect 81452 16574 81480 50322
rect 82832 16574 82860 76502
rect 107580 75886 107608 91287
rect 108946 91216 109002 91225
rect 108304 91180 108356 91186
rect 108946 91151 109002 91160
rect 109590 91216 109646 91225
rect 109590 91151 109646 91160
rect 108304 91122 108356 91128
rect 108316 81394 108344 91122
rect 108304 81388 108356 81394
rect 108304 81330 108356 81336
rect 108960 79966 108988 91151
rect 109604 86766 109632 91151
rect 109592 86760 109644 86766
rect 109592 86702 109644 86708
rect 110156 82618 110184 93191
rect 115480 92472 115532 92478
rect 115478 92440 115480 92449
rect 115532 92440 115534 92449
rect 115478 92375 115534 92384
rect 116766 92440 116822 92449
rect 116766 92375 116822 92384
rect 120538 92440 120594 92449
rect 122852 92410 122880 94454
rect 129384 94042 129412 94687
rect 151648 94110 151676 94687
rect 161478 94480 161534 94489
rect 161478 94415 161534 94424
rect 151636 94104 151688 94110
rect 151636 94046 151688 94052
rect 129372 94036 129424 94042
rect 129372 93978 129424 93984
rect 133142 93664 133198 93673
rect 133142 93599 133198 93608
rect 133156 93430 133184 93599
rect 133144 93424 133196 93430
rect 133144 93366 133196 93372
rect 125506 92440 125562 92449
rect 120538 92375 120594 92384
rect 122840 92404 122892 92410
rect 116780 92342 116808 92375
rect 116768 92336 116820 92342
rect 110326 92304 110382 92313
rect 116768 92278 116820 92284
rect 110326 92239 110382 92248
rect 110340 90846 110368 92239
rect 115386 91760 115442 91769
rect 115386 91695 115442 91704
rect 111430 91352 111486 91361
rect 111430 91287 111486 91296
rect 114374 91352 114430 91361
rect 114374 91287 114430 91296
rect 111246 91216 111302 91225
rect 111246 91151 111302 91160
rect 110328 90840 110380 90846
rect 110328 90782 110380 90788
rect 111260 88126 111288 91151
rect 111248 88120 111300 88126
rect 111248 88062 111300 88068
rect 111444 85474 111472 91287
rect 112350 91216 112406 91225
rect 112350 91151 112406 91160
rect 112364 86698 112392 91151
rect 114388 88233 114416 91287
rect 114466 91216 114522 91225
rect 114466 91151 114522 91160
rect 114374 88224 114430 88233
rect 114374 88159 114430 88168
rect 112352 86692 112404 86698
rect 112352 86634 112404 86640
rect 111432 85468 111484 85474
rect 111432 85410 111484 85416
rect 110144 82612 110196 82618
rect 110144 82554 110196 82560
rect 108948 79960 109000 79966
rect 108948 79902 109000 79908
rect 114480 79830 114508 91151
rect 115400 89418 115428 91695
rect 115846 91216 115902 91225
rect 115846 91151 115902 91160
rect 117134 91216 117190 91225
rect 117134 91151 117190 91160
rect 118606 91216 118662 91225
rect 118606 91151 118662 91160
rect 119986 91216 120042 91225
rect 119986 91151 120042 91160
rect 115388 89412 115440 89418
rect 115388 89354 115440 89360
rect 115860 80034 115888 91151
rect 117148 88058 117176 91151
rect 117136 88052 117188 88058
rect 117136 87994 117188 88000
rect 118620 84114 118648 91151
rect 118608 84108 118660 84114
rect 118608 84050 118660 84056
rect 115848 80028 115900 80034
rect 115848 79970 115900 79976
rect 114468 79824 114520 79830
rect 114468 79766 114520 79772
rect 120000 78470 120028 91151
rect 120552 90982 120580 92375
rect 125506 92375 125562 92384
rect 125966 92440 126022 92449
rect 125966 92375 125968 92384
rect 122840 92346 122892 92352
rect 122838 91488 122894 91497
rect 122838 91423 122894 91432
rect 122746 91352 122802 91361
rect 122746 91287 122802 91296
rect 122654 91216 122710 91225
rect 122654 91151 122710 91160
rect 120540 90976 120592 90982
rect 120540 90918 120592 90924
rect 122668 83842 122696 91151
rect 122656 83836 122708 83842
rect 122656 83778 122708 83784
rect 122760 82822 122788 91287
rect 122852 85270 122880 91423
rect 123482 91216 123538 91225
rect 123482 91151 123538 91160
rect 124126 91216 124182 91225
rect 124126 91151 124182 91160
rect 125414 91216 125470 91225
rect 125414 91151 125470 91160
rect 123496 87990 123524 91151
rect 123484 87984 123536 87990
rect 123484 87926 123536 87932
rect 124140 86630 124168 91151
rect 124128 86624 124180 86630
rect 124128 86566 124180 86572
rect 122840 85264 122892 85270
rect 122840 85206 122892 85212
rect 122748 82816 122800 82822
rect 122748 82758 122800 82764
rect 125428 82482 125456 91151
rect 125520 90778 125548 92375
rect 126020 92375 126022 92384
rect 130750 92440 130806 92449
rect 130750 92375 130806 92384
rect 151726 92440 151782 92449
rect 151726 92375 151782 92384
rect 152094 92440 152150 92449
rect 152094 92375 152150 92384
rect 125968 92346 126020 92352
rect 130764 92206 130792 92375
rect 151740 92274 151768 92375
rect 151728 92268 151780 92274
rect 151728 92210 151780 92216
rect 130752 92200 130804 92206
rect 130752 92142 130804 92148
rect 136454 92168 136510 92177
rect 152108 92138 152136 92375
rect 136454 92103 136510 92112
rect 152096 92132 152148 92138
rect 126702 91760 126758 91769
rect 126702 91695 126758 91704
rect 126518 91216 126574 91225
rect 126518 91151 126574 91160
rect 125508 90772 125560 90778
rect 125508 90714 125560 90720
rect 126532 88194 126560 91151
rect 126716 89729 126744 91695
rect 128266 91216 128322 91225
rect 128266 91151 128322 91160
rect 132406 91216 132462 91225
rect 132406 91151 132462 91160
rect 134614 91216 134670 91225
rect 134614 91151 134670 91160
rect 126702 89720 126758 89729
rect 126702 89655 126758 89664
rect 126520 88188 126572 88194
rect 126520 88130 126572 88136
rect 125416 82476 125468 82482
rect 125416 82418 125468 82424
rect 128280 81258 128308 91151
rect 129004 91112 129056 91118
rect 129004 91054 129056 91060
rect 128268 81252 128320 81258
rect 128268 81194 128320 81200
rect 129016 78606 129044 91054
rect 132420 85202 132448 91151
rect 134628 86834 134656 91151
rect 136468 90710 136496 92103
rect 152096 92074 152148 92080
rect 161492 91633 161520 94415
rect 161478 91624 161534 91633
rect 161478 91559 161534 91568
rect 151266 91488 151322 91497
rect 151266 91423 151322 91432
rect 136456 90704 136508 90710
rect 136456 90646 136508 90652
rect 151280 89350 151308 91423
rect 151268 89344 151320 89350
rect 151268 89286 151320 89292
rect 134616 86828 134668 86834
rect 134616 86770 134668 86776
rect 132408 85196 132460 85202
rect 132408 85138 132460 85144
rect 129004 78600 129056 78606
rect 129004 78542 129056 78548
rect 119988 78464 120040 78470
rect 119988 78406 120040 78412
rect 124220 76628 124272 76634
rect 124220 76570 124272 76576
rect 107568 75880 107620 75886
rect 107568 75822 107620 75828
rect 115940 75268 115992 75274
rect 115940 75210 115992 75216
rect 93860 73908 93912 73914
rect 93860 73850 93912 73856
rect 85580 57248 85632 57254
rect 85580 57190 85632 57196
rect 84200 43512 84252 43518
rect 84200 43454 84252 43460
rect 77404 16546 78168 16574
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 77312 6886 77432 6914
rect 77404 480 77432 6886
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 43454
rect 85592 6914 85620 57190
rect 86960 53168 87012 53174
rect 86960 53110 87012 53116
rect 85672 21480 85724 21486
rect 85672 21422 85724 21428
rect 85684 16574 85712 21422
rect 86972 16574 87000 53110
rect 91100 51808 91152 51814
rect 91100 51750 91152 51756
rect 88340 47592 88392 47598
rect 88340 47534 88392 47540
rect 88352 16574 88380 47534
rect 89720 18624 89772 18630
rect 89720 18566 89772 18572
rect 89732 16574 89760 18566
rect 91112 16574 91140 51750
rect 92480 36644 92532 36650
rect 92480 36586 92532 36592
rect 85684 16546 86448 16574
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 85592 6886 85712 6914
rect 85684 480 85712 6886
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 36586
rect 93872 6914 93900 73850
rect 103520 71120 103572 71126
rect 103520 71062 103572 71068
rect 98000 61396 98052 61402
rect 98000 61338 98052 61344
rect 93952 44940 94004 44946
rect 93952 44882 94004 44888
rect 93964 16574 93992 44882
rect 95240 43444 95292 43450
rect 95240 43386 95292 43392
rect 95252 16574 95280 43386
rect 96620 26988 96672 26994
rect 96620 26930 96672 26936
rect 96632 16574 96660 26930
rect 98012 16574 98040 61338
rect 102140 49088 102192 49094
rect 102140 49030 102192 49036
rect 99380 38004 99432 38010
rect 99380 37946 99432 37952
rect 99392 16574 99420 37946
rect 100760 22840 100812 22846
rect 100760 22782 100812 22788
rect 93964 16546 94728 16574
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 93872 6886 93992 6914
rect 93964 480 93992 6886
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 22782
rect 102152 16574 102180 49030
rect 103532 16574 103560 71062
rect 110420 68400 110472 68406
rect 110420 68342 110472 68348
rect 104900 50448 104952 50454
rect 104900 50390 104952 50396
rect 104912 16574 104940 50390
rect 106280 33856 106332 33862
rect 106280 33798 106332 33804
rect 106292 16574 106320 33798
rect 107660 24200 107712 24206
rect 107660 24142 107712 24148
rect 107672 16574 107700 24142
rect 102152 16546 102272 16574
rect 103532 16546 104112 16574
rect 104912 16546 105768 16574
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 102244 480 102272 16546
rect 103336 7676 103388 7682
rect 103336 7618 103388 7624
rect 103348 480 103376 7618
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105740 480 105768 16546
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 110432 3602 110460 68342
rect 114560 66972 114612 66978
rect 114560 66914 114612 66920
rect 114572 16574 114600 66914
rect 115952 16574 115980 75210
rect 118700 72548 118752 72554
rect 118700 72490 118752 72496
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 110512 3664 110564 3670
rect 110512 3606 110564 3612
rect 112812 3664 112864 3670
rect 112812 3606 112864 3612
rect 110420 3596 110472 3602
rect 110420 3538 110472 3544
rect 109316 2100 109368 2106
rect 109316 2042 109368 2048
rect 109328 480 109356 2042
rect 110524 480 110552 3606
rect 111616 3596 111668 3602
rect 111616 3538 111668 3544
rect 111628 480 111656 3538
rect 112824 480 112852 3606
rect 114008 2168 114060 2174
rect 114008 2110 114060 2116
rect 114020 480 114048 2110
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 117320 10396 117372 10402
rect 117320 10338 117372 10344
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 10338
rect 118712 3398 118740 72490
rect 121460 65612 121512 65618
rect 121460 65554 121512 65560
rect 118792 25628 118844 25634
rect 118792 25570 118844 25576
rect 118700 3392 118752 3398
rect 118700 3334 118752 3340
rect 118804 480 118832 25570
rect 121472 16574 121500 65554
rect 122840 46232 122892 46238
rect 122840 46174 122892 46180
rect 122852 16574 122880 46174
rect 124232 16574 124260 76570
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 124232 16546 124720 16574
rect 120632 11824 120684 11830
rect 120632 11766 120684 11772
rect 119896 3392 119948 3398
rect 119896 3334 119948 3340
rect 119908 480 119936 3334
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 11766
rect 122300 480 122328 16546
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124692 480 124720 16546
rect 164896 3738 164924 95095
rect 164988 93158 165016 97990
rect 166276 94042 166304 143550
rect 167644 140820 167696 140826
rect 167644 140762 167696 140768
rect 166906 115832 166962 115841
rect 166906 115767 166962 115776
rect 166540 99476 166592 99482
rect 166540 99418 166592 99424
rect 166356 99408 166408 99414
rect 166356 99350 166408 99356
rect 166264 94036 166316 94042
rect 166264 93978 166316 93984
rect 164976 93152 165028 93158
rect 164976 93094 165028 93100
rect 166368 82754 166396 99350
rect 166448 98116 166500 98122
rect 166448 98058 166500 98064
rect 166460 84046 166488 98058
rect 166552 86902 166580 99418
rect 166920 98025 166948 115767
rect 166906 98016 166962 98025
rect 166906 97951 166962 97960
rect 166540 86896 166592 86902
rect 166540 86838 166592 86844
rect 166448 84040 166500 84046
rect 166448 83982 166500 83988
rect 166356 82748 166408 82754
rect 166356 82690 166408 82696
rect 167656 82482 167684 140762
rect 167748 90710 167776 147630
rect 173164 145036 173216 145042
rect 173164 144978 173216 144984
rect 169024 144968 169076 144974
rect 169024 144910 169076 144916
rect 167828 133952 167880 133958
rect 167828 133894 167880 133900
rect 167736 90704 167788 90710
rect 167736 90646 167788 90652
rect 167840 88126 167868 133894
rect 167920 118720 167972 118726
rect 167920 118662 167972 118668
rect 167828 88120 167880 88126
rect 167828 88062 167880 88068
rect 167932 86698 167960 118662
rect 168012 111784 168064 111790
rect 168010 111752 168012 111761
rect 168064 111752 168066 111761
rect 168010 111687 168066 111696
rect 168104 110424 168156 110430
rect 168104 110366 168156 110372
rect 168116 110129 168144 110366
rect 168102 110120 168158 110129
rect 168102 110055 168158 110064
rect 168012 108996 168064 109002
rect 168012 108938 168064 108944
rect 168024 108769 168052 108938
rect 168010 108760 168066 108769
rect 168010 108695 168066 108704
rect 169036 92206 169064 144910
rect 171784 139460 171836 139466
rect 171784 139402 171836 139408
rect 170404 138032 170456 138038
rect 170404 137974 170456 137980
rect 169116 125656 169168 125662
rect 169116 125598 169168 125604
rect 169024 92200 169076 92206
rect 169024 92142 169076 92148
rect 169128 90778 169156 125598
rect 169208 111852 169260 111858
rect 169208 111794 169260 111800
rect 169116 90772 169168 90778
rect 169116 90714 169168 90720
rect 167920 86692 167972 86698
rect 167920 86634 167972 86640
rect 169220 85338 169248 111794
rect 169300 106344 169352 106350
rect 169300 106286 169352 106292
rect 169208 85332 169260 85338
rect 169208 85274 169260 85280
rect 167644 82476 167696 82482
rect 167644 82418 167696 82424
rect 169312 81326 169340 106286
rect 170416 93362 170444 137974
rect 170496 135312 170548 135318
rect 170496 135254 170548 135260
rect 170508 93974 170536 135254
rect 170588 124228 170640 124234
rect 170588 124170 170640 124176
rect 170496 93968 170548 93974
rect 170496 93910 170548 93916
rect 170404 93356 170456 93362
rect 170404 93298 170456 93304
rect 170600 86630 170628 124170
rect 170680 120148 170732 120154
rect 170680 120090 170732 120096
rect 170692 88058 170720 120090
rect 170680 88052 170732 88058
rect 170680 87994 170732 88000
rect 170588 86624 170640 86630
rect 170588 86566 170640 86572
rect 171796 83842 171824 139402
rect 171968 137284 172020 137290
rect 171968 137226 172020 137232
rect 171876 129804 171928 129810
rect 171876 129746 171928 129752
rect 171784 83836 171836 83842
rect 171784 83778 171836 83784
rect 171888 82550 171916 129746
rect 171980 111790 172008 137226
rect 172060 118788 172112 118794
rect 172060 118730 172112 118736
rect 171968 111784 172020 111790
rect 171968 111726 172020 111732
rect 171968 103556 172020 103562
rect 171968 103498 172020 103504
rect 171980 91050 172008 103498
rect 172072 93906 172100 118730
rect 172060 93900 172112 93906
rect 172060 93842 172112 93848
rect 171968 91044 172020 91050
rect 171968 90986 172020 90992
rect 173176 85202 173204 144978
rect 173268 92138 173296 151030
rect 175924 150476 175976 150482
rect 175924 150418 175976 150424
rect 174544 146328 174596 146334
rect 174544 146270 174596 146276
rect 173348 132524 173400 132530
rect 173348 132466 173400 132472
rect 173256 92132 173308 92138
rect 173256 92074 173308 92080
rect 173164 85196 173216 85202
rect 173164 85138 173216 85144
rect 171876 82544 171928 82550
rect 171876 82486 171928 82492
rect 169300 81320 169352 81326
rect 169300 81262 169352 81268
rect 173360 81190 173388 132466
rect 173440 110492 173492 110498
rect 173440 110434 173492 110440
rect 173452 82686 173480 110434
rect 174556 93430 174584 146270
rect 174728 117972 174780 117978
rect 174728 117914 174780 117920
rect 174636 109064 174688 109070
rect 174636 109006 174688 109012
rect 174544 93424 174596 93430
rect 174544 93366 174596 93372
rect 174648 83978 174676 109006
rect 174740 92342 174768 117914
rect 175936 110430 175964 150418
rect 176108 116000 176160 116006
rect 176108 115942 176160 115948
rect 176016 114572 176068 114578
rect 176016 114514 176068 114520
rect 175924 110424 175976 110430
rect 175924 110366 175976 110372
rect 174728 92336 174780 92342
rect 174728 92278 174780 92284
rect 174636 83972 174688 83978
rect 174636 83914 174688 83920
rect 173440 82680 173492 82686
rect 173440 82622 173492 82628
rect 173348 81184 173400 81190
rect 173348 81126 173400 81132
rect 176028 75886 176056 114514
rect 176120 90846 176148 115942
rect 177316 95169 177344 294199
rect 178684 292732 178736 292738
rect 178684 292674 178736 292680
rect 178696 177313 178724 292674
rect 180064 269136 180116 269142
rect 180064 269078 180116 269084
rect 180076 184346 180104 269078
rect 184204 224324 184256 224330
rect 184204 224266 184256 224272
rect 180064 184340 180116 184346
rect 180064 184282 180116 184288
rect 178682 177304 178738 177313
rect 178682 177239 178738 177248
rect 178684 153264 178736 153270
rect 178684 153206 178736 153212
rect 177580 151836 177632 151842
rect 177580 151778 177632 151784
rect 177396 140888 177448 140894
rect 177396 140830 177448 140836
rect 177302 95160 177358 95169
rect 177302 95095 177358 95104
rect 176108 90840 176160 90846
rect 176108 90782 176160 90788
rect 177304 90364 177356 90370
rect 177304 90306 177356 90312
rect 176016 75880 176068 75886
rect 176016 75822 176068 75828
rect 125876 3732 125928 3738
rect 125876 3674 125928 3680
rect 164884 3732 164936 3738
rect 164884 3674 164936 3680
rect 125888 480 125916 3674
rect 177316 3534 177344 90306
rect 177408 87990 177436 140830
rect 177488 134020 177540 134026
rect 177488 133962 177540 133968
rect 177396 87984 177448 87990
rect 177396 87926 177448 87932
rect 177500 86766 177528 133962
rect 177592 109002 177620 151778
rect 177580 108996 177632 109002
rect 177580 108938 177632 108944
rect 177672 107704 177724 107710
rect 177672 107646 177724 107652
rect 177488 86760 177540 86766
rect 177488 86702 177540 86708
rect 177684 79898 177712 107646
rect 178696 94110 178724 153206
rect 178776 128376 178828 128382
rect 178776 128318 178828 128324
rect 178684 94104 178736 94110
rect 178684 94046 178736 94052
rect 177672 79892 177724 79898
rect 177672 79834 177724 79840
rect 178788 78538 178816 128318
rect 180064 124296 180116 124302
rect 180064 124238 180116 124244
rect 178868 118856 178920 118862
rect 178868 118798 178920 118804
rect 178880 89418 178908 118798
rect 178868 89412 178920 89418
rect 178868 89354 178920 89360
rect 180076 85270 180104 124238
rect 182824 121508 182876 121514
rect 182824 121450 182876 121456
rect 181444 117360 181496 117366
rect 181444 117302 181496 117308
rect 180156 114640 180208 114646
rect 180156 114582 180208 114588
rect 180064 85264 180116 85270
rect 180064 85206 180116 85212
rect 180168 83910 180196 114582
rect 180156 83904 180208 83910
rect 180156 83846 180208 83852
rect 181456 82618 181484 117302
rect 181444 82612 181496 82618
rect 181444 82554 181496 82560
rect 178776 78532 178828 78538
rect 178776 78474 178828 78480
rect 182836 78470 182864 121450
rect 182824 78464 182876 78470
rect 182824 78406 182876 78412
rect 184216 60722 184244 224266
rect 186976 182986 187004 298386
rect 198004 298376 198056 298382
rect 198004 298318 198056 298324
rect 188342 294128 188398 294137
rect 188342 294063 188398 294072
rect 186964 182980 187016 182986
rect 186964 182922 187016 182928
rect 186962 176896 187018 176905
rect 186962 176831 187018 176840
rect 186976 158642 187004 176831
rect 186964 158636 187016 158642
rect 186964 158578 187016 158584
rect 186964 116068 187016 116074
rect 186964 116010 187016 116016
rect 186976 93226 187004 116010
rect 188356 93770 188384 294063
rect 195244 281648 195296 281654
rect 195244 281590 195296 281596
rect 191196 233912 191248 233918
rect 191196 233854 191248 233860
rect 191104 205080 191156 205086
rect 191104 205022 191156 205028
rect 189724 131164 189776 131170
rect 189724 131106 189776 131112
rect 188344 93764 188396 93770
rect 188344 93706 188396 93712
rect 186964 93220 187016 93226
rect 186964 93162 187016 93168
rect 189736 90914 189764 131106
rect 191116 93702 191144 205022
rect 191208 180266 191236 233854
rect 191196 180260 191248 180266
rect 191196 180202 191248 180208
rect 195256 177342 195284 281590
rect 196624 238128 196676 238134
rect 196624 238070 196676 238076
rect 195244 177336 195296 177342
rect 195244 177278 195296 177284
rect 195336 176724 195388 176730
rect 195336 176666 195388 176672
rect 195348 161362 195376 176666
rect 195336 161356 195388 161362
rect 195336 161298 195388 161304
rect 195244 135380 195296 135386
rect 195244 135322 195296 135328
rect 191196 125724 191248 125730
rect 191196 125666 191248 125672
rect 191104 93696 191156 93702
rect 191104 93638 191156 93644
rect 189724 90908 189776 90914
rect 189724 90850 189776 90856
rect 191208 88194 191236 125666
rect 192484 110560 192536 110566
rect 192484 110502 192536 110508
rect 192496 89486 192524 110502
rect 192484 89480 192536 89486
rect 192484 89422 192536 89428
rect 191196 88188 191248 88194
rect 191196 88130 191248 88136
rect 195256 79830 195284 135322
rect 195336 122868 195388 122874
rect 195336 122810 195388 122816
rect 195348 93294 195376 122810
rect 196636 95198 196664 238070
rect 198016 185609 198044 298318
rect 198002 185600 198058 185609
rect 198002 185535 198058 185544
rect 202156 181626 202184 299610
rect 204904 295588 204956 295594
rect 204904 295530 204956 295536
rect 202144 181620 202196 181626
rect 202144 181562 202196 181568
rect 204916 178770 204944 295530
rect 206296 187066 206324 299678
rect 209044 249824 209096 249830
rect 209044 249766 209096 249772
rect 206284 187060 206336 187066
rect 206284 187002 206336 187008
rect 209056 178906 209084 249766
rect 213196 183054 213224 302398
rect 214576 233238 214604 699654
rect 235184 698970 235212 703520
rect 235172 698964 235224 698970
rect 235172 698906 235224 698912
rect 267660 697678 267688 703520
rect 266360 697672 266412 697678
rect 266360 697614 266412 697620
rect 267648 697672 267700 697678
rect 267648 697614 267700 697620
rect 233884 305108 233936 305114
rect 233884 305050 233936 305056
rect 224224 302388 224276 302394
rect 224224 302330 224276 302336
rect 220084 300960 220136 300966
rect 220084 300902 220136 300908
rect 215944 297016 215996 297022
rect 215944 296958 215996 296964
rect 214656 236700 214708 236706
rect 214656 236642 214708 236648
rect 214564 233232 214616 233238
rect 214564 233174 214616 233180
rect 214668 188562 214696 236642
rect 214656 188556 214708 188562
rect 214656 188498 214708 188504
rect 214564 187740 214616 187746
rect 214564 187682 214616 187688
rect 213184 183048 213236 183054
rect 213184 182990 213236 182996
rect 213276 182232 213328 182238
rect 213276 182174 213328 182180
rect 211804 179444 211856 179450
rect 211804 179386 211856 179392
rect 209044 178900 209096 178906
rect 209044 178842 209096 178848
rect 204904 178764 204956 178770
rect 204904 178706 204956 178712
rect 209044 175976 209096 175982
rect 209044 175918 209096 175924
rect 209056 157282 209084 175918
rect 211816 171018 211844 179386
rect 211896 176792 211948 176798
rect 211896 176734 211948 176740
rect 211804 171012 211856 171018
rect 211804 170954 211856 170960
rect 211908 169658 211936 176734
rect 212264 176112 212316 176118
rect 212264 176054 212316 176060
rect 212276 172514 212304 176054
rect 212264 172508 212316 172514
rect 212264 172450 212316 172456
rect 213288 172417 213316 182174
rect 213920 176860 213972 176866
rect 213920 176802 213972 176808
rect 213932 176225 213960 176802
rect 213918 176216 213974 176225
rect 213918 176151 213974 176160
rect 213920 175228 213972 175234
rect 213920 175170 213972 175176
rect 213932 175137 213960 175170
rect 213918 175128 213974 175137
rect 213918 175063 213974 175072
rect 214576 174729 214604 187682
rect 214656 186380 214708 186386
rect 214656 186322 214708 186328
rect 214562 174720 214618 174729
rect 214562 174655 214618 174664
rect 214668 174570 214696 186322
rect 215956 178838 215984 296958
rect 216036 202224 216088 202230
rect 216036 202166 216088 202172
rect 215944 178832 215996 178838
rect 215944 178774 215996 178780
rect 214748 176044 214800 176050
rect 214748 175986 214800 175992
rect 214012 174548 214064 174554
rect 214012 174490 214064 174496
rect 214392 174542 214696 174570
rect 213920 173868 213972 173874
rect 213920 173810 213972 173816
rect 213932 173777 213960 173810
rect 213918 173768 213974 173777
rect 213918 173703 213974 173712
rect 214024 173369 214052 174490
rect 214010 173360 214066 173369
rect 214010 173295 214066 173304
rect 213920 172508 213972 172514
rect 213920 172450 213972 172456
rect 213274 172408 213330 172417
rect 213274 172343 213330 172352
rect 213932 172009 213960 172450
rect 213918 172000 213974 172009
rect 213918 171935 213974 171944
rect 213920 171080 213972 171086
rect 213920 171022 213972 171028
rect 213932 170785 213960 171022
rect 213918 170776 213974 170785
rect 213918 170711 213974 170720
rect 214392 169810 214420 174542
rect 214656 173188 214708 173194
rect 214656 173130 214708 173136
rect 214472 171148 214524 171154
rect 214524 171106 214604 171134
rect 214472 171090 214524 171096
rect 214472 171012 214524 171018
rect 214472 170954 214524 170960
rect 214484 170921 214512 170954
rect 214470 170912 214526 170921
rect 214470 170847 214526 170856
rect 214392 169782 214512 169810
rect 213920 169720 213972 169726
rect 213920 169662 213972 169668
rect 214010 169688 214066 169697
rect 211896 169652 211948 169658
rect 211896 169594 211948 169600
rect 213932 169425 213960 169662
rect 214010 169623 214012 169632
rect 214064 169623 214066 169632
rect 214012 169594 214064 169600
rect 213918 169416 213974 169425
rect 213918 169351 213974 169360
rect 213920 168360 213972 168366
rect 213920 168302 213972 168308
rect 213932 168065 213960 168302
rect 214012 168292 214064 168298
rect 214012 168234 214064 168240
rect 213918 168056 213974 168065
rect 213918 167991 213974 168000
rect 214024 167929 214052 168234
rect 214010 167920 214066 167929
rect 214010 167855 214066 167864
rect 213920 167000 213972 167006
rect 213920 166942 213972 166948
rect 213932 166161 213960 166942
rect 214484 166705 214512 169782
rect 214470 166696 214526 166705
rect 214470 166631 214526 166640
rect 213918 166152 213974 166161
rect 213918 166087 213974 166096
rect 213920 165572 213972 165578
rect 213920 165514 213972 165520
rect 213932 165345 213960 165514
rect 214012 165504 214064 165510
rect 214012 165446 214064 165452
rect 213918 165336 213974 165345
rect 213918 165271 213974 165280
rect 214024 164801 214052 165446
rect 214010 164792 214066 164801
rect 214010 164727 214066 164736
rect 214012 164212 214064 164218
rect 214012 164154 214064 164160
rect 213920 164144 213972 164150
rect 213918 164112 213920 164121
rect 213972 164112 213974 164121
rect 213918 164047 213974 164056
rect 214024 163441 214052 164154
rect 214010 163432 214066 163441
rect 214010 163367 214066 163376
rect 213920 162852 213972 162858
rect 213920 162794 213972 162800
rect 213932 161537 213960 162794
rect 213918 161528 213974 161537
rect 213918 161463 213974 161472
rect 214012 161424 214064 161430
rect 214012 161366 214064 161372
rect 213920 161356 213972 161362
rect 213920 161298 213972 161304
rect 213932 161265 213960 161298
rect 213918 161256 213974 161265
rect 213918 161191 213974 161200
rect 214024 160857 214052 161366
rect 214010 160848 214066 160857
rect 214010 160783 214066 160792
rect 213920 160064 213972 160070
rect 213918 160032 213920 160041
rect 213972 160032 213974 160041
rect 213918 159967 213974 159976
rect 213920 158704 213972 158710
rect 213918 158672 213920 158681
rect 213972 158672 213974 158681
rect 213918 158607 213974 158616
rect 214012 158636 214064 158642
rect 214012 158578 214064 158584
rect 214024 158137 214052 158578
rect 214010 158128 214066 158137
rect 214010 158063 214066 158072
rect 214012 157344 214064 157350
rect 213918 157312 213974 157321
rect 209044 157276 209096 157282
rect 214012 157286 214064 157292
rect 213918 157247 213920 157256
rect 209044 157218 209096 157224
rect 213972 157247 213974 157256
rect 213920 157218 213972 157224
rect 214024 156913 214052 157286
rect 214010 156904 214066 156913
rect 214010 156839 214066 156848
rect 213920 155916 213972 155922
rect 213920 155858 213972 155864
rect 213932 155553 213960 155858
rect 213918 155544 213974 155553
rect 213918 155479 213974 155488
rect 214010 153912 214066 153921
rect 214010 153847 214066 153856
rect 213918 153504 213974 153513
rect 213918 153439 213974 153448
rect 198004 153332 198056 153338
rect 198004 153274 198056 153280
rect 196716 132592 196768 132598
rect 196716 132534 196768 132540
rect 196624 95192 196676 95198
rect 196624 95134 196676 95140
rect 195336 93288 195388 93294
rect 195336 93230 195388 93236
rect 196728 79966 196756 132534
rect 198016 92274 198044 153274
rect 213932 153270 213960 153439
rect 214024 153338 214052 153847
rect 214012 153332 214064 153338
rect 214012 153274 214064 153280
rect 213920 153264 213972 153270
rect 213920 153206 213972 153212
rect 213182 152688 213238 152697
rect 213182 152623 213238 152632
rect 210424 146396 210476 146402
rect 210424 146338 210476 146344
rect 202144 143676 202196 143682
rect 202144 143618 202196 143624
rect 199384 129872 199436 129878
rect 199384 129814 199436 129820
rect 198096 113212 198148 113218
rect 198096 113154 198148 113160
rect 198004 92268 198056 92274
rect 198004 92210 198056 92216
rect 198108 85406 198136 113154
rect 198188 95260 198240 95266
rect 198188 95202 198240 95208
rect 198096 85400 198148 85406
rect 198096 85342 198148 85348
rect 196716 79960 196768 79966
rect 196716 79902 196768 79908
rect 195244 79824 195296 79830
rect 195244 79766 195296 79772
rect 198200 77246 198228 95202
rect 199396 94489 199424 129814
rect 199476 104916 199528 104922
rect 199476 104858 199528 104864
rect 199382 94480 199438 94489
rect 199382 94415 199438 94424
rect 199488 89622 199516 104858
rect 199476 89616 199528 89622
rect 199476 89558 199528 89564
rect 202156 81258 202184 143618
rect 206376 142180 206428 142186
rect 206376 142122 206428 142128
rect 204904 136672 204956 136678
rect 204904 136614 204956 136620
rect 202236 121576 202288 121582
rect 202236 121518 202288 121524
rect 202248 84114 202276 121518
rect 204916 92478 204944 136614
rect 204996 111920 205048 111926
rect 204996 111862 205048 111868
rect 204904 92472 204956 92478
rect 204904 92414 204956 92420
rect 205008 86970 205036 111862
rect 206388 92410 206416 142122
rect 209044 139528 209096 139534
rect 209044 139470 209096 139476
rect 207664 131232 207716 131238
rect 207664 131174 207716 131180
rect 206376 92404 206428 92410
rect 206376 92346 206428 92352
rect 206284 91792 206336 91798
rect 206284 91734 206336 91740
rect 204996 86964 205048 86970
rect 204996 86906 205048 86912
rect 202236 84108 202288 84114
rect 202236 84050 202288 84056
rect 202144 81252 202196 81258
rect 202144 81194 202196 81200
rect 198188 77240 198240 77246
rect 198188 77182 198240 77188
rect 184204 60716 184256 60722
rect 184204 60658 184256 60664
rect 206296 3670 206324 91734
rect 207676 84182 207704 131174
rect 207756 104984 207808 104990
rect 207756 104926 207808 104932
rect 207768 94897 207796 104926
rect 207754 94888 207810 94897
rect 207754 94823 207810 94832
rect 209056 90982 209084 139470
rect 209136 109132 209188 109138
rect 209136 109074 209188 109080
rect 209044 90976 209096 90982
rect 209044 90918 209096 90924
rect 207664 84176 207716 84182
rect 207664 84118 207716 84124
rect 209148 78674 209176 109074
rect 210436 86834 210464 146338
rect 211804 123412 211856 123418
rect 211804 123354 211856 123360
rect 210608 103896 210660 103902
rect 210608 103838 210660 103844
rect 210516 96688 210568 96694
rect 210516 96630 210568 96636
rect 210424 86828 210476 86834
rect 210424 86770 210476 86776
rect 210528 85542 210556 96630
rect 210620 93838 210648 103838
rect 210608 93832 210660 93838
rect 210608 93774 210660 93780
rect 210516 85536 210568 85542
rect 210516 85478 210568 85484
rect 211816 82822 211844 123354
rect 211896 113280 211948 113286
rect 211896 113222 211948 113228
rect 211908 89554 211936 113222
rect 211896 89548 211948 89554
rect 211896 89490 211948 89496
rect 213196 89350 213224 152623
rect 214378 152144 214434 152153
rect 214378 152079 214434 152088
rect 213918 152008 213974 152017
rect 213918 151943 213974 151952
rect 213932 151842 213960 151943
rect 213920 151836 213972 151842
rect 213920 151778 213972 151784
rect 214392 151094 214420 152079
rect 214380 151088 214432 151094
rect 214380 151030 214432 151036
rect 214010 150920 214066 150929
rect 214010 150855 214066 150864
rect 214024 150482 214052 150855
rect 214012 150476 214064 150482
rect 214012 150418 214064 150424
rect 213920 150408 213972 150414
rect 213920 150350 213972 150356
rect 213932 150113 213960 150350
rect 213918 150104 213974 150113
rect 213918 150039 213974 150048
rect 214576 149569 214604 171106
rect 214668 159497 214696 173130
rect 214760 166977 214788 175986
rect 214746 166968 214802 166977
rect 214746 166903 214802 166912
rect 214654 159488 214710 159497
rect 214654 159423 214710 159432
rect 214654 150784 214710 150793
rect 214654 150719 214710 150728
rect 214562 149560 214618 149569
rect 214562 149495 214618 149504
rect 213920 149048 213972 149054
rect 213920 148990 213972 148996
rect 213932 148753 213960 148990
rect 213918 148744 213974 148753
rect 213918 148679 213974 148688
rect 213918 148064 213974 148073
rect 213918 147999 213974 148008
rect 213932 147694 213960 147999
rect 213920 147688 213972 147694
rect 213920 147630 213972 147636
rect 214010 146704 214066 146713
rect 214010 146639 214066 146648
rect 213918 146432 213974 146441
rect 214024 146402 214052 146639
rect 213918 146367 213974 146376
rect 214012 146396 214064 146402
rect 213932 146334 213960 146367
rect 214012 146338 214064 146344
rect 213920 146328 213972 146334
rect 213920 146270 213972 146276
rect 214010 145344 214066 145353
rect 214010 145279 214066 145288
rect 214024 145042 214052 145279
rect 214012 145036 214064 145042
rect 214012 144978 214064 144984
rect 213920 144968 213972 144974
rect 213918 144936 213920 144945
rect 213972 144936 213974 144945
rect 213918 144871 213974 144880
rect 214010 143984 214066 143993
rect 214010 143919 214066 143928
rect 213920 143676 213972 143682
rect 213920 143618 213972 143624
rect 213932 143585 213960 143618
rect 214024 143614 214052 143919
rect 214012 143608 214064 143614
rect 213918 143576 213974 143585
rect 214012 143550 214064 143556
rect 213918 143511 213974 143520
rect 213918 142216 213974 142225
rect 213918 142151 213920 142160
rect 213972 142151 213974 142160
rect 214668 142154 214696 150719
rect 213920 142122 213972 142128
rect 214576 142126 214696 142154
rect 214010 141400 214066 141409
rect 214010 141335 214066 141344
rect 213918 140992 213974 141001
rect 213918 140927 213974 140936
rect 213932 140894 213960 140927
rect 213920 140888 213972 140894
rect 213920 140830 213972 140836
rect 214024 140826 214052 141335
rect 214012 140820 214064 140826
rect 214012 140762 214064 140768
rect 214010 140040 214066 140049
rect 214010 139975 214066 139984
rect 213918 139632 213974 139641
rect 213918 139567 213974 139576
rect 213932 139534 213960 139567
rect 213920 139528 213972 139534
rect 213920 139470 213972 139476
rect 214024 139466 214052 139975
rect 214012 139460 214064 139466
rect 214012 139402 214064 139408
rect 214470 138816 214526 138825
rect 214470 138751 214526 138760
rect 213918 138136 213974 138145
rect 213918 138071 213974 138080
rect 213932 138038 213960 138071
rect 213920 138032 213972 138038
rect 213920 137974 213972 137980
rect 213918 136776 213974 136785
rect 213918 136711 213974 136720
rect 213932 136678 213960 136711
rect 213920 136672 213972 136678
rect 213920 136614 213972 136620
rect 214010 135688 214066 135697
rect 214010 135623 214066 135632
rect 213918 135416 213974 135425
rect 214024 135386 214052 135623
rect 213918 135351 213974 135360
rect 214012 135380 214064 135386
rect 213932 135318 213960 135351
rect 214012 135322 214064 135328
rect 213920 135312 213972 135318
rect 213920 135254 213972 135260
rect 214010 134328 214066 134337
rect 214010 134263 214066 134272
rect 213918 134056 213974 134065
rect 213918 133991 213920 134000
rect 213972 133991 213974 134000
rect 213920 133962 213972 133968
rect 214024 133958 214052 134263
rect 214012 133952 214064 133958
rect 214012 133894 214064 133900
rect 214010 132832 214066 132841
rect 214010 132767 214066 132776
rect 214024 132598 214052 132767
rect 214012 132592 214064 132598
rect 213918 132560 213974 132569
rect 214012 132534 214064 132540
rect 213918 132495 213920 132504
rect 213972 132495 213974 132504
rect 213920 132466 213972 132472
rect 214484 132494 214512 138751
rect 214576 137290 214604 142126
rect 214654 137456 214710 137465
rect 214654 137391 214710 137400
rect 214564 137284 214616 137290
rect 214564 137226 214616 137232
rect 214668 132494 214696 137391
rect 214484 132466 214604 132494
rect 214668 132466 214788 132494
rect 214010 131472 214066 131481
rect 214010 131407 214066 131416
rect 213920 131232 213972 131238
rect 213918 131200 213920 131209
rect 213972 131200 213974 131209
rect 214024 131170 214052 131407
rect 213918 131135 213974 131144
rect 214012 131164 214064 131170
rect 214012 131106 214064 131112
rect 214010 130112 214066 130121
rect 214010 130047 214066 130056
rect 214024 129878 214052 130047
rect 214012 129872 214064 129878
rect 213918 129840 213974 129849
rect 214012 129814 214064 129820
rect 213918 129775 213920 129784
rect 213972 129775 213974 129784
rect 213920 129746 213972 129752
rect 213918 128888 213974 128897
rect 213918 128823 213974 128832
rect 213932 128382 213960 128823
rect 213920 128376 213972 128382
rect 213920 128318 213972 128324
rect 213458 127528 213514 127537
rect 213458 127463 213514 127472
rect 213472 127129 213500 127463
rect 213458 127120 213514 127129
rect 213458 127055 213514 127064
rect 214010 126168 214066 126177
rect 214010 126103 214066 126112
rect 213918 125760 213974 125769
rect 214024 125730 214052 126103
rect 213918 125695 213974 125704
rect 214012 125724 214064 125730
rect 213932 125662 213960 125695
rect 214012 125666 214064 125672
rect 213920 125656 213972 125662
rect 213920 125598 213972 125604
rect 214010 124808 214066 124817
rect 214010 124743 214066 124752
rect 213918 124400 213974 124409
rect 213918 124335 213974 124344
rect 213932 124302 213960 124335
rect 213920 124296 213972 124302
rect 213920 124238 213972 124244
rect 214024 124234 214052 124743
rect 214012 124228 214064 124234
rect 214012 124170 214064 124176
rect 213918 123584 213974 123593
rect 213918 123519 213974 123528
rect 213932 123418 213960 123519
rect 213920 123412 213972 123418
rect 213920 123354 213972 123360
rect 213918 122904 213974 122913
rect 213918 122839 213920 122848
rect 213972 122839 213974 122848
rect 213920 122810 213972 122816
rect 214010 122224 214066 122233
rect 214010 122159 214066 122168
rect 213918 121816 213974 121825
rect 213918 121751 213974 121760
rect 213932 121582 213960 121751
rect 213920 121576 213972 121582
rect 213920 121518 213972 121524
rect 214024 121514 214052 122159
rect 214012 121508 214064 121514
rect 214012 121450 214064 121456
rect 213918 120864 213974 120873
rect 213918 120799 213974 120808
rect 213274 120184 213330 120193
rect 213932 120154 213960 120799
rect 213274 120119 213330 120128
rect 213920 120148 213972 120154
rect 213184 89344 213236 89350
rect 213184 89286 213236 89292
rect 211804 82816 211856 82822
rect 211804 82758 211856 82764
rect 213288 80034 213316 120119
rect 213920 120090 213972 120096
rect 214010 119640 214066 119649
rect 214010 119575 214066 119584
rect 213918 118960 213974 118969
rect 213918 118895 213974 118904
rect 213932 118726 213960 118895
rect 214024 118862 214052 119575
rect 214102 119096 214158 119105
rect 214102 119031 214158 119040
rect 214012 118856 214064 118862
rect 214012 118798 214064 118804
rect 214116 118794 214144 119031
rect 214104 118788 214156 118794
rect 214104 118730 214156 118736
rect 213920 118720 213972 118726
rect 213920 118662 213972 118668
rect 213366 117600 213422 117609
rect 213366 117535 213422 117544
rect 213380 85474 213408 117535
rect 213920 117360 213972 117366
rect 213918 117328 213920 117337
rect 213972 117328 213974 117337
rect 213918 117263 213974 117272
rect 214010 116240 214066 116249
rect 214010 116175 214066 116184
rect 213920 116068 213972 116074
rect 213920 116010 213972 116016
rect 213932 115977 213960 116010
rect 214024 116006 214052 116175
rect 214012 116000 214064 116006
rect 213918 115968 213974 115977
rect 214012 115942 214064 115948
rect 213918 115903 213974 115912
rect 214010 115016 214066 115025
rect 214010 114951 214066 114960
rect 213920 114640 213972 114646
rect 213918 114608 213920 114617
rect 213972 114608 213974 114617
rect 214024 114578 214052 114951
rect 213918 114543 213974 114552
rect 214012 114572 214064 114578
rect 214012 114514 214064 114520
rect 213918 113656 213974 113665
rect 213918 113591 213974 113600
rect 213932 113218 213960 113591
rect 214012 113280 214064 113286
rect 214010 113248 214012 113257
rect 214064 113248 214066 113257
rect 213920 113212 213972 113218
rect 214010 113183 214066 113192
rect 213920 113154 213972 113160
rect 214010 112296 214066 112305
rect 214010 112231 214066 112240
rect 214024 111926 214052 112231
rect 214012 111920 214064 111926
rect 213918 111888 213974 111897
rect 214012 111862 214064 111868
rect 213918 111823 213920 111832
rect 213972 111823 213974 111832
rect 213920 111794 213972 111800
rect 214010 110936 214066 110945
rect 214010 110871 214066 110880
rect 214024 110566 214052 110871
rect 214012 110560 214064 110566
rect 213918 110528 213974 110537
rect 214012 110502 214064 110508
rect 213918 110463 213920 110472
rect 213972 110463 213974 110472
rect 213920 110434 213972 110440
rect 214010 109712 214066 109721
rect 214010 109647 214066 109656
rect 213918 109304 213974 109313
rect 213918 109239 213974 109248
rect 213932 109070 213960 109239
rect 214024 109138 214052 109647
rect 214012 109132 214064 109138
rect 214012 109074 214064 109080
rect 213920 109064 213972 109070
rect 213920 109006 213972 109012
rect 213918 107944 213974 107953
rect 213918 107879 213974 107888
rect 213932 107710 213960 107879
rect 213920 107704 213972 107710
rect 213920 107646 213972 107652
rect 213918 106992 213974 107001
rect 213918 106927 213974 106936
rect 213932 106350 213960 106927
rect 213920 106344 213972 106350
rect 213920 106286 213972 106292
rect 214010 105768 214066 105777
rect 214010 105703 214066 105712
rect 213918 105360 213974 105369
rect 213918 105295 213974 105304
rect 213932 104990 213960 105295
rect 213920 104984 213972 104990
rect 213920 104926 213972 104932
rect 214024 104922 214052 105703
rect 214012 104916 214064 104922
rect 214012 104858 214064 104864
rect 213918 104000 213974 104009
rect 213918 103935 213974 103944
rect 213932 103902 213960 103935
rect 213920 103896 213972 103902
rect 213920 103838 213972 103844
rect 213918 103728 213974 103737
rect 213918 103663 213974 103672
rect 213932 103562 213960 103663
rect 213920 103556 213972 103562
rect 214576 103514 214604 132466
rect 214760 117978 214788 132466
rect 214748 117972 214800 117978
rect 214748 117914 214800 117920
rect 214838 108352 214894 108361
rect 214838 108287 214894 108296
rect 214654 106312 214710 106321
rect 214654 106247 214710 106256
rect 213920 103498 213972 103504
rect 214484 103486 214604 103514
rect 214010 99784 214066 99793
rect 214010 99719 214066 99728
rect 213918 99512 213974 99521
rect 213918 99447 213920 99456
rect 213972 99447 213974 99456
rect 213920 99418 213972 99424
rect 214024 99414 214052 99719
rect 214012 99408 214064 99414
rect 214012 99350 214064 99356
rect 214010 98424 214066 98433
rect 214010 98359 214066 98368
rect 214024 98122 214052 98359
rect 214012 98116 214064 98122
rect 214012 98058 214064 98064
rect 213920 98048 213972 98054
rect 213918 98016 213920 98025
rect 213972 98016 213974 98025
rect 213918 97951 213974 97960
rect 214484 97209 214512 103486
rect 214562 101144 214618 101153
rect 214562 101079 214618 101088
rect 214470 97200 214526 97209
rect 214470 97135 214526 97144
rect 213918 97064 213974 97073
rect 213918 96999 213974 97008
rect 213932 96694 213960 96999
rect 213920 96688 213972 96694
rect 213920 96630 213972 96636
rect 213918 95840 213974 95849
rect 213918 95775 213974 95784
rect 213932 95266 213960 95775
rect 213920 95260 213972 95266
rect 213920 95202 213972 95208
rect 214576 88262 214604 101079
rect 214564 88256 214616 88262
rect 214564 88198 214616 88204
rect 213368 85468 213420 85474
rect 213368 85410 213420 85416
rect 214668 81394 214696 106247
rect 214852 94518 214880 108287
rect 214930 96656 214986 96665
rect 214930 96591 214986 96600
rect 214840 94512 214892 94518
rect 214840 94454 214892 94460
rect 214944 88330 214972 96591
rect 216048 93838 216076 202166
rect 220096 175953 220124 300902
rect 222844 240236 222896 240242
rect 222844 240178 222896 240184
rect 222856 180334 222884 240178
rect 222844 180328 222896 180334
rect 222844 180270 222896 180276
rect 224236 176089 224264 302330
rect 226984 298308 227036 298314
rect 226984 298250 227036 298256
rect 226996 177449 227024 298250
rect 231124 278860 231176 278866
rect 231124 278802 231176 278808
rect 228364 273284 228416 273290
rect 228364 273226 228416 273232
rect 228376 180402 228404 273226
rect 228364 180396 228416 180402
rect 228364 180338 228416 180344
rect 231136 178974 231164 278802
rect 232504 256760 232556 256766
rect 232504 256702 232556 256708
rect 231124 178968 231176 178974
rect 231124 178910 231176 178916
rect 232516 177585 232544 256702
rect 232502 177576 232558 177585
rect 232502 177511 232558 177520
rect 226982 177440 227038 177449
rect 226982 177375 227038 177384
rect 224222 176080 224278 176089
rect 224222 176015 224278 176024
rect 233896 175982 233924 305050
rect 244924 303748 244976 303754
rect 244924 303690 244976 303696
rect 242164 281580 242216 281586
rect 242164 281522 242216 281528
rect 238024 243568 238076 243574
rect 238024 243510 238076 243516
rect 233976 213240 234028 213246
rect 233976 213182 234028 213188
rect 233988 177410 234016 213182
rect 238036 180470 238064 243510
rect 238116 211880 238168 211886
rect 238116 211822 238168 211828
rect 238128 183122 238156 211822
rect 240784 210452 240836 210458
rect 240784 210394 240836 210400
rect 238116 183116 238168 183122
rect 238116 183058 238168 183064
rect 238024 180464 238076 180470
rect 238024 180406 238076 180412
rect 233976 177404 234028 177410
rect 233976 177346 234028 177352
rect 240796 176050 240824 210394
rect 242176 178022 242204 281522
rect 244936 183190 244964 303690
rect 252560 295520 252612 295526
rect 252560 295462 252612 295468
rect 250444 284368 250496 284374
rect 250444 284310 250496 284316
rect 246304 259480 246356 259486
rect 246304 259422 246356 259428
rect 245016 217456 245068 217462
rect 245016 217398 245068 217404
rect 244924 183184 244976 183190
rect 244924 183126 244976 183132
rect 245028 178809 245056 217398
rect 245014 178800 245070 178809
rect 245014 178735 245070 178744
rect 242164 178016 242216 178022
rect 242164 177958 242216 177964
rect 246316 177478 246344 259422
rect 250456 199646 250484 284310
rect 251180 232552 251232 232558
rect 251180 232494 251232 232500
rect 250444 199640 250496 199646
rect 250444 199582 250496 199588
rect 249800 196648 249852 196654
rect 249800 196590 249852 196596
rect 246948 181620 247000 181626
rect 246948 181562 247000 181568
rect 246304 177472 246356 177478
rect 246304 177414 246356 177420
rect 240784 176044 240836 176050
rect 240784 175986 240836 175992
rect 233884 175976 233936 175982
rect 220082 175944 220138 175953
rect 233884 175918 233936 175924
rect 220082 175879 220138 175888
rect 246960 175817 246988 181562
rect 249064 178968 249116 178974
rect 249064 178910 249116 178916
rect 246946 175808 247002 175817
rect 246946 175743 247002 175752
rect 249076 172786 249104 178910
rect 249248 178900 249300 178906
rect 249248 178842 249300 178848
rect 249156 178016 249208 178022
rect 249156 177958 249208 177964
rect 249168 174729 249196 177958
rect 249260 175273 249288 178842
rect 249246 175264 249302 175273
rect 249246 175199 249302 175208
rect 249154 174720 249210 174729
rect 249154 174655 249210 174664
rect 249154 172800 249210 172809
rect 249076 172758 249154 172786
rect 249154 172735 249210 172744
rect 217322 155408 217378 155417
rect 217322 155343 217378 155352
rect 217336 154737 217364 155343
rect 217322 154728 217378 154737
rect 217322 154663 217378 154672
rect 249812 150793 249840 196590
rect 249892 191412 249944 191418
rect 249892 191354 249944 191360
rect 249904 165753 249932 191354
rect 249984 175976 250036 175982
rect 249984 175918 250036 175924
rect 249890 165744 249946 165753
rect 249890 165679 249946 165688
rect 249996 161474 250024 175918
rect 249904 161446 250024 161474
rect 249904 158273 249932 161446
rect 251192 158817 251220 232494
rect 251272 194132 251324 194138
rect 251272 194074 251324 194080
rect 251178 158808 251234 158817
rect 251178 158743 251234 158752
rect 249890 158264 249946 158273
rect 249890 158199 249946 158208
rect 250442 155272 250498 155281
rect 250442 155207 250498 155216
rect 249798 150784 249854 150793
rect 249798 150719 249854 150728
rect 250456 143721 250484 155207
rect 251284 151814 251312 194074
rect 251364 177336 251416 177342
rect 251364 177278 251416 177284
rect 251376 160177 251404 177278
rect 252466 173768 252522 173777
rect 252466 173703 252522 173712
rect 252480 172582 252508 173703
rect 252468 172576 252520 172582
rect 252468 172518 252520 172524
rect 252374 172408 252430 172417
rect 252374 172343 252430 172352
rect 252468 172372 252520 172378
rect 252388 171426 252416 172343
rect 252468 172314 252520 172320
rect 252480 171465 252508 172314
rect 252466 171456 252522 171465
rect 252376 171420 252428 171426
rect 252466 171391 252522 171400
rect 252376 171362 252428 171368
rect 252468 170808 252520 170814
rect 252468 170750 252520 170756
rect 252480 170241 252508 170750
rect 252466 170232 252522 170241
rect 252466 170167 252522 170176
rect 252466 170096 252522 170105
rect 252466 170031 252522 170040
rect 252480 169862 252508 170031
rect 252468 169856 252520 169862
rect 252468 169798 252520 169804
rect 252376 169720 252428 169726
rect 252376 169662 252428 169668
rect 252284 169652 252336 169658
rect 252284 169594 252336 169600
rect 252296 168609 252324 169594
rect 252388 169153 252416 169662
rect 252466 169552 252522 169561
rect 252466 169487 252522 169496
rect 252374 169144 252430 169153
rect 252374 169079 252430 169088
rect 252480 168978 252508 169487
rect 252468 168972 252520 168978
rect 252468 168914 252520 168920
rect 252282 168600 252338 168609
rect 252282 168535 252338 168544
rect 252376 168360 252428 168366
rect 252376 168302 252428 168308
rect 252284 168292 252336 168298
rect 252284 168234 252336 168240
rect 252296 167657 252324 168234
rect 252282 167648 252338 167657
rect 252282 167583 252338 167592
rect 252388 167249 252416 168302
rect 252466 168192 252522 168201
rect 252466 168127 252522 168136
rect 252480 167890 252508 168127
rect 252468 167884 252520 167890
rect 252468 167826 252520 167832
rect 252374 167240 252430 167249
rect 252374 167175 252430 167184
rect 252466 166696 252522 166705
rect 252466 166631 252522 166640
rect 252374 166288 252430 166297
rect 252480 166258 252508 166631
rect 252374 166223 252430 166232
rect 252468 166252 252520 166258
rect 252388 165782 252416 166223
rect 252468 166194 252520 166200
rect 252376 165776 252428 165782
rect 252376 165718 252428 165724
rect 252376 165572 252428 165578
rect 252376 165514 252428 165520
rect 252388 164801 252416 165514
rect 252468 165504 252520 165510
rect 252468 165446 252520 165452
rect 252480 165345 252508 165446
rect 252466 165336 252522 165345
rect 252466 165271 252522 165280
rect 252374 164792 252430 164801
rect 252374 164727 252430 164736
rect 252468 164212 252520 164218
rect 252468 164154 252520 164160
rect 251456 164144 251508 164150
rect 251456 164086 251508 164092
rect 251468 163033 251496 164086
rect 252480 163985 252508 164154
rect 252466 163976 252522 163985
rect 252466 163911 252522 163920
rect 251454 163024 251510 163033
rect 251454 162959 251510 162968
rect 252376 162852 252428 162858
rect 252376 162794 252428 162800
rect 252284 162784 252336 162790
rect 252284 162726 252336 162732
rect 252296 161537 252324 162726
rect 252388 162081 252416 162794
rect 252468 162716 252520 162722
rect 252468 162658 252520 162664
rect 252480 162489 252508 162658
rect 252466 162480 252522 162489
rect 252466 162415 252522 162424
rect 252374 162072 252430 162081
rect 252374 162007 252430 162016
rect 252282 161528 252338 161537
rect 252282 161463 252338 161472
rect 252468 160812 252520 160818
rect 252468 160754 252520 160760
rect 252480 160585 252508 160754
rect 252466 160576 252522 160585
rect 252466 160511 252522 160520
rect 251362 160168 251418 160177
rect 251362 160103 251418 160112
rect 252468 160064 252520 160070
rect 252468 160006 252520 160012
rect 252008 159996 252060 160002
rect 252008 159938 252060 159944
rect 252020 159225 252048 159938
rect 252480 159633 252508 160006
rect 252466 159624 252522 159633
rect 252466 159559 252522 159568
rect 252006 159216 252062 159225
rect 252006 159151 252062 159160
rect 252468 157344 252520 157350
rect 252466 157312 252468 157321
rect 252520 157312 252522 157321
rect 252376 157276 252428 157282
rect 252466 157247 252522 157256
rect 252376 157218 252428 157224
rect 252388 156369 252416 157218
rect 252468 157208 252520 157214
rect 252468 157150 252520 157156
rect 252480 156913 252508 157150
rect 252466 156904 252522 156913
rect 252466 156839 252522 156848
rect 252374 156360 252430 156369
rect 252374 156295 252430 156304
rect 252466 155952 252522 155961
rect 252376 155916 252428 155922
rect 252466 155887 252522 155896
rect 252376 155858 252428 155864
rect 251456 155780 251508 155786
rect 251456 155722 251508 155728
rect 251468 155417 251496 155722
rect 251454 155408 251510 155417
rect 251454 155343 251510 155352
rect 252388 155009 252416 155858
rect 252480 155854 252508 155887
rect 252468 155848 252520 155854
rect 252468 155790 252520 155796
rect 252374 155000 252430 155009
rect 252374 154935 252430 154944
rect 252376 154556 252428 154562
rect 252376 154498 252428 154504
rect 252284 154420 252336 154426
rect 252284 154362 252336 154368
rect 252296 152153 252324 154362
rect 252388 154057 252416 154498
rect 252468 154488 252520 154494
rect 252466 154456 252468 154465
rect 252520 154456 252522 154465
rect 252466 154391 252522 154400
rect 252374 154048 252430 154057
rect 252374 153983 252430 153992
rect 252468 153128 252520 153134
rect 252466 153096 252468 153105
rect 252520 153096 252522 153105
rect 252466 153031 252522 153040
rect 252572 152697 252600 295462
rect 255412 294160 255464 294166
rect 255412 294102 255464 294108
rect 255320 289944 255372 289950
rect 255320 289886 255372 289892
rect 252652 268388 252704 268394
rect 252652 268330 252704 268336
rect 252664 171873 252692 268330
rect 253940 263628 253992 263634
rect 253940 263570 253992 263576
rect 252744 221536 252796 221542
rect 252744 221478 252796 221484
rect 252650 171864 252706 171873
rect 252650 171799 252706 171808
rect 252756 164393 252784 221478
rect 252836 181484 252888 181490
rect 252836 181426 252888 181432
rect 252742 164384 252798 164393
rect 252742 164319 252798 164328
rect 252558 152688 252614 152697
rect 252558 152623 252614 152632
rect 252282 152144 252338 152153
rect 252282 152079 252338 152088
rect 251284 151786 251404 151814
rect 251272 147552 251324 147558
rect 251272 147494 251324 147500
rect 251284 146985 251312 147494
rect 251270 146976 251326 146985
rect 251270 146911 251326 146920
rect 250442 143712 250498 143721
rect 250442 143647 250498 143656
rect 251376 140865 251404 151786
rect 252468 151768 252520 151774
rect 252466 151736 252468 151745
rect 252520 151736 252522 151745
rect 252466 151671 252522 151680
rect 252008 151496 252060 151502
rect 252008 151438 252060 151444
rect 252020 151201 252048 151438
rect 252006 151192 252062 151201
rect 252006 151127 252062 151136
rect 252468 150408 252520 150414
rect 252468 150350 252520 150356
rect 252376 150340 252428 150346
rect 252376 150282 252428 150288
rect 252284 150272 252336 150278
rect 252282 150240 252284 150249
rect 252336 150240 252338 150249
rect 252282 150175 252338 150184
rect 252388 149297 252416 150282
rect 252480 149841 252508 150350
rect 252466 149832 252522 149841
rect 252466 149767 252522 149776
rect 252374 149288 252430 149297
rect 252374 149223 252430 149232
rect 252468 149048 252520 149054
rect 252468 148990 252520 148996
rect 252376 148980 252428 148986
rect 252376 148922 252428 148928
rect 252388 147937 252416 148922
rect 252480 148345 252508 148990
rect 252848 148889 252876 181426
rect 253952 164150 253980 263570
rect 254124 222896 254176 222902
rect 254124 222838 254176 222844
rect 254032 214668 254084 214674
rect 254032 214610 254084 214616
rect 253940 164144 253992 164150
rect 253940 164086 253992 164092
rect 253204 161492 253256 161498
rect 253204 161434 253256 161440
rect 252834 148880 252890 148889
rect 252834 148815 252890 148824
rect 252466 148336 252522 148345
rect 252466 148271 252522 148280
rect 252374 147928 252430 147937
rect 252374 147863 252430 147872
rect 252468 147620 252520 147626
rect 252468 147562 252520 147568
rect 252480 146577 252508 147562
rect 252466 146568 252522 146577
rect 252466 146503 252522 146512
rect 252190 146296 252246 146305
rect 252190 146231 252246 146240
rect 252284 146260 252336 146266
rect 252008 145580 252060 145586
rect 252008 145522 252060 145528
rect 251916 142860 251968 142866
rect 251916 142802 251968 142808
rect 251362 140856 251418 140865
rect 251362 140791 251418 140800
rect 250444 138032 250496 138038
rect 250444 137974 250496 137980
rect 216218 102504 216274 102513
rect 216218 102439 216274 102448
rect 216126 100872 216182 100881
rect 216126 100807 216182 100816
rect 216036 93832 216088 93838
rect 216036 93774 216088 93780
rect 215944 89004 215996 89010
rect 215944 88946 215996 88952
rect 214932 88324 214984 88330
rect 214932 88266 214984 88272
rect 214656 81388 214708 81394
rect 214656 81330 214708 81336
rect 213276 80028 213328 80034
rect 213276 79970 213328 79976
rect 209136 78668 209188 78674
rect 209136 78610 209188 78616
rect 206284 3664 206336 3670
rect 206284 3606 206336 3612
rect 215956 3602 215984 88946
rect 216140 78606 216168 100807
rect 216232 89690 216260 102439
rect 249154 96656 249210 96665
rect 249154 96591 249210 96600
rect 249064 95260 249116 95266
rect 249064 95202 249116 95208
rect 238024 91860 238076 91866
rect 238024 91802 238076 91808
rect 216220 89684 216272 89690
rect 216220 89626 216272 89632
rect 216128 78600 216180 78606
rect 216128 78542 216180 78548
rect 215944 3596 215996 3602
rect 215944 3538 215996 3544
rect 238036 3534 238064 91802
rect 249076 60042 249104 95202
rect 249064 60036 249116 60042
rect 249064 59978 249116 59984
rect 249168 46918 249196 96591
rect 249156 46912 249208 46918
rect 249156 46854 249208 46860
rect 250456 11830 250484 137974
rect 251824 137352 251876 137358
rect 251824 137294 251876 137300
rect 251836 122834 251864 137294
rect 251928 126313 251956 142802
rect 252020 136241 252048 145522
rect 252204 142769 252232 146231
rect 252284 146202 252336 146208
rect 252296 145081 252324 146202
rect 252468 146192 252520 146198
rect 252468 146134 252520 146140
rect 252376 146124 252428 146130
rect 252376 146066 252428 146072
rect 252388 145625 252416 146066
rect 252480 146033 252508 146134
rect 252466 146024 252522 146033
rect 252466 145959 252522 145968
rect 252374 145616 252430 145625
rect 252374 145551 252430 145560
rect 252282 145072 252338 145081
rect 252282 145007 252338 145016
rect 252468 144900 252520 144906
rect 252468 144842 252520 144848
rect 252480 144129 252508 144842
rect 252466 144120 252522 144129
rect 252466 144055 252522 144064
rect 252376 143540 252428 143546
rect 252376 143482 252428 143488
rect 252190 142760 252246 142769
rect 252190 142695 252246 142704
rect 252388 142225 252416 143482
rect 252468 143472 252520 143478
rect 252468 143414 252520 143420
rect 252480 143177 252508 143414
rect 252466 143168 252522 143177
rect 252466 143103 252522 143112
rect 252374 142216 252430 142225
rect 252374 142151 252430 142160
rect 252468 142112 252520 142118
rect 252468 142054 252520 142060
rect 252480 141409 252508 142054
rect 252466 141400 252522 141409
rect 252466 141335 252522 141344
rect 252468 140752 252520 140758
rect 252468 140694 252520 140700
rect 252376 140684 252428 140690
rect 252376 140626 252428 140632
rect 252388 139505 252416 140626
rect 252480 139913 252508 140694
rect 252466 139904 252522 139913
rect 252466 139839 252522 139848
rect 252374 139496 252430 139505
rect 252374 139431 252430 139440
rect 252284 139392 252336 139398
rect 252284 139334 252336 139340
rect 252192 138712 252244 138718
rect 252192 138654 252244 138660
rect 252006 136232 252062 136241
rect 252006 136167 252062 136176
rect 252204 132841 252232 138654
rect 252296 138553 252324 139334
rect 252282 138544 252338 138553
rect 252282 138479 252338 138488
rect 252374 138000 252430 138009
rect 252284 137964 252336 137970
rect 252374 137935 252430 137944
rect 252284 137906 252336 137912
rect 252296 137057 252324 137906
rect 252388 137902 252416 137935
rect 252376 137896 252428 137902
rect 252376 137838 252428 137844
rect 252468 137828 252520 137834
rect 252468 137770 252520 137776
rect 252480 137601 252508 137770
rect 252466 137592 252522 137601
rect 252466 137527 252522 137536
rect 252282 137048 252338 137057
rect 252282 136983 252338 136992
rect 252466 136640 252522 136649
rect 252284 136604 252336 136610
rect 252466 136575 252522 136584
rect 252284 136546 252336 136552
rect 252296 135697 252324 136546
rect 252480 136542 252508 136575
rect 252468 136536 252520 136542
rect 252468 136478 252520 136484
rect 252376 136468 252428 136474
rect 252376 136410 252428 136416
rect 252282 135688 252338 135697
rect 252282 135623 252338 135632
rect 252388 135289 252416 136410
rect 252374 135280 252430 135289
rect 252374 135215 252430 135224
rect 252468 135244 252520 135250
rect 252468 135186 252520 135192
rect 252376 135176 252428 135182
rect 252376 135118 252428 135124
rect 252388 134337 252416 135118
rect 252480 134745 252508 135186
rect 252466 134736 252522 134745
rect 252466 134671 252522 134680
rect 252374 134328 252430 134337
rect 252374 134263 252430 134272
rect 252376 133884 252428 133890
rect 252376 133826 252428 133832
rect 252388 133385 252416 133826
rect 252468 133816 252520 133822
rect 252466 133784 252468 133793
rect 252520 133784 252522 133793
rect 252466 133719 252522 133728
rect 252374 133376 252430 133385
rect 252374 133311 252430 133320
rect 252190 132832 252246 132841
rect 252190 132767 252246 132776
rect 252284 132456 252336 132462
rect 252284 132398 252336 132404
rect 252374 132424 252430 132433
rect 252296 131481 252324 132398
rect 252374 132359 252430 132368
rect 252468 132388 252520 132394
rect 252388 131578 252416 132359
rect 252468 132330 252520 132336
rect 252480 131889 252508 132330
rect 252466 131880 252522 131889
rect 252466 131815 252522 131824
rect 252376 131572 252428 131578
rect 252376 131514 252428 131520
rect 252282 131472 252338 131481
rect 252282 131407 252338 131416
rect 252284 131096 252336 131102
rect 252284 131038 252336 131044
rect 252296 130121 252324 131038
rect 252468 131028 252520 131034
rect 252468 130970 252520 130976
rect 252480 130529 252508 130970
rect 252466 130520 252522 130529
rect 252466 130455 252522 130464
rect 252376 130416 252428 130422
rect 252376 130358 252428 130364
rect 252282 130112 252338 130121
rect 252282 130047 252338 130056
rect 252284 129668 252336 129674
rect 252284 129610 252336 129616
rect 252008 129056 252060 129062
rect 252008 128998 252060 129004
rect 251914 126304 251970 126313
rect 251914 126239 251970 126248
rect 251652 122806 251864 122834
rect 251652 117337 251680 122806
rect 251916 120760 251968 120766
rect 251916 120702 251968 120708
rect 251638 117328 251694 117337
rect 251638 117263 251694 117272
rect 251928 110809 251956 120702
rect 252020 116929 252048 128998
rect 252296 128625 252324 129610
rect 252388 129577 252416 130358
rect 252468 129736 252520 129742
rect 252468 129678 252520 129684
rect 252374 129568 252430 129577
rect 252374 129503 252430 129512
rect 252480 129169 252508 129678
rect 252466 129160 252522 129169
rect 252466 129095 252522 129104
rect 252282 128616 252338 128625
rect 252282 128551 252338 128560
rect 252376 128308 252428 128314
rect 252376 128250 252428 128256
rect 252388 127673 252416 128250
rect 252468 128240 252520 128246
rect 252466 128208 252468 128217
rect 252520 128208 252522 128217
rect 252466 128143 252522 128152
rect 252374 127664 252430 127673
rect 252374 127599 252430 127608
rect 252468 127492 252520 127498
rect 252468 127434 252520 127440
rect 252480 127265 252508 127434
rect 252466 127256 252522 127265
rect 252466 127191 252522 127200
rect 252468 126948 252520 126954
rect 252468 126890 252520 126896
rect 252480 126721 252508 126890
rect 252466 126712 252522 126721
rect 252376 126676 252428 126682
rect 252466 126647 252522 126656
rect 252376 126618 252428 126624
rect 252192 126268 252244 126274
rect 252192 126210 252244 126216
rect 252204 124409 252232 126210
rect 252388 125769 252416 126618
rect 252374 125760 252430 125769
rect 252374 125695 252430 125704
rect 252468 125588 252520 125594
rect 252468 125530 252520 125536
rect 252376 125520 252428 125526
rect 252376 125462 252428 125468
rect 252388 125361 252416 125462
rect 252374 125352 252430 125361
rect 252374 125287 252430 125296
rect 252284 124908 252336 124914
rect 252284 124850 252336 124856
rect 252190 124400 252246 124409
rect 252190 124335 252246 124344
rect 252296 124001 252324 124850
rect 252480 124817 252508 125530
rect 252466 124808 252522 124817
rect 252466 124743 252522 124752
rect 252468 124160 252520 124166
rect 252468 124102 252520 124108
rect 252376 124092 252428 124098
rect 252376 124034 252428 124040
rect 252282 123992 252338 124001
rect 252282 123927 252338 123936
rect 252284 123480 252336 123486
rect 252284 123422 252336 123428
rect 252296 120193 252324 123422
rect 252388 123049 252416 124034
rect 252480 123457 252508 124102
rect 252466 123448 252522 123457
rect 252466 123383 252522 123392
rect 252374 123040 252430 123049
rect 252374 122975 252430 122984
rect 252376 122732 252428 122738
rect 252376 122674 252428 122680
rect 252388 121553 252416 122674
rect 252468 122664 252520 122670
rect 252468 122606 252520 122612
rect 252480 122505 252508 122606
rect 252466 122496 252522 122505
rect 252466 122431 252522 122440
rect 253216 122097 253244 161434
rect 254044 147558 254072 214610
rect 254136 155786 254164 222838
rect 254216 198076 254268 198082
rect 254216 198018 254268 198024
rect 254124 155780 254176 155786
rect 254124 155722 254176 155728
rect 254228 151502 254256 198018
rect 255332 160002 255360 289886
rect 255424 168298 255452 294102
rect 262220 280288 262272 280294
rect 262220 280230 262272 280236
rect 255504 274712 255556 274718
rect 255504 274654 255556 274660
rect 255412 168292 255464 168298
rect 255412 168234 255464 168240
rect 255320 159996 255372 160002
rect 255320 159938 255372 159944
rect 255516 154426 255544 274654
rect 259736 220176 259788 220182
rect 259736 220118 259788 220124
rect 258080 199572 258132 199578
rect 258080 199514 258132 199520
rect 256792 183184 256844 183190
rect 256792 183126 256844 183132
rect 255596 180260 255648 180266
rect 255596 180202 255648 180208
rect 255504 154420 255556 154426
rect 255504 154362 255556 154368
rect 254216 151496 254268 151502
rect 254216 151438 254268 151444
rect 254584 150476 254636 150482
rect 254584 150418 254636 150424
rect 254032 147552 254084 147558
rect 254032 147494 254084 147500
rect 253296 143608 253348 143614
rect 253296 143550 253348 143556
rect 253202 122088 253258 122097
rect 253202 122023 253258 122032
rect 252374 121544 252430 121553
rect 252374 121479 252430 121488
rect 252376 121440 252428 121446
rect 252376 121382 252428 121388
rect 252388 120601 252416 121382
rect 252466 121136 252522 121145
rect 252466 121071 252522 121080
rect 252480 120698 252508 121071
rect 252468 120692 252520 120698
rect 252468 120634 252520 120640
rect 252374 120592 252430 120601
rect 252374 120527 252430 120536
rect 252282 120184 252338 120193
rect 252282 120119 252338 120128
rect 252376 120080 252428 120086
rect 252376 120022 252428 120028
rect 252388 118833 252416 120022
rect 252468 120012 252520 120018
rect 252468 119954 252520 119960
rect 252480 119649 252508 119954
rect 252466 119640 252522 119649
rect 252466 119575 252522 119584
rect 252468 119468 252520 119474
rect 252468 119410 252520 119416
rect 252480 119241 252508 119410
rect 252466 119232 252522 119241
rect 252466 119167 252522 119176
rect 252374 118824 252430 118833
rect 252374 118759 252430 118768
rect 252468 118652 252520 118658
rect 252468 118594 252520 118600
rect 252376 118584 252428 118590
rect 252376 118526 252428 118532
rect 252284 117972 252336 117978
rect 252284 117914 252336 117920
rect 252006 116920 252062 116929
rect 252006 116855 252062 116864
rect 252100 116612 252152 116618
rect 252100 116554 252152 116560
rect 252008 112464 252060 112470
rect 252008 112406 252060 112412
rect 251914 110800 251970 110809
rect 251914 110735 251970 110744
rect 251640 110288 251692 110294
rect 251640 110230 251692 110236
rect 251652 109857 251680 110230
rect 251638 109848 251694 109857
rect 251638 109783 251694 109792
rect 251272 104168 251324 104174
rect 251272 104110 251324 104116
rect 251180 103352 251232 103358
rect 251180 103294 251232 103300
rect 251192 103193 251220 103294
rect 251178 103184 251234 103193
rect 251178 103119 251234 103128
rect 251284 98569 251312 104110
rect 252020 103737 252048 112406
rect 252112 108905 252140 116554
rect 252296 115433 252324 117914
rect 252388 117881 252416 118526
rect 252480 118289 252508 118594
rect 252466 118280 252522 118289
rect 252466 118215 252522 118224
rect 252374 117872 252430 117881
rect 252374 117807 252430 117816
rect 252468 117292 252520 117298
rect 252468 117234 252520 117240
rect 252480 116385 252508 117234
rect 252466 116376 252522 116385
rect 252466 116311 252522 116320
rect 252468 116136 252520 116142
rect 252468 116078 252520 116084
rect 252480 115977 252508 116078
rect 252466 115968 252522 115977
rect 252376 115932 252428 115938
rect 252466 115903 252522 115912
rect 252376 115874 252428 115880
rect 252282 115424 252338 115433
rect 252282 115359 252338 115368
rect 252284 115252 252336 115258
rect 252284 115194 252336 115200
rect 252296 113529 252324 115194
rect 252388 115025 252416 115874
rect 252374 115016 252430 115025
rect 252374 114951 252430 114960
rect 252468 114504 252520 114510
rect 252466 114472 252468 114481
rect 252520 114472 252522 114481
rect 252376 114436 252428 114442
rect 252466 114407 252522 114416
rect 252376 114378 252428 114384
rect 252388 114073 252416 114378
rect 252374 114064 252430 114073
rect 252374 113999 252430 114008
rect 252282 113520 252338 113529
rect 252282 113455 252338 113464
rect 252468 113144 252520 113150
rect 252468 113086 252520 113092
rect 252480 112169 252508 113086
rect 252466 112160 252522 112169
rect 252466 112095 252522 112104
rect 253204 111852 253256 111858
rect 253204 111794 253256 111800
rect 252468 111784 252520 111790
rect 252374 111752 252430 111761
rect 252468 111726 252520 111732
rect 252374 111687 252376 111696
rect 252428 111687 252430 111696
rect 252376 111658 252428 111664
rect 252480 111217 252508 111726
rect 252466 111208 252522 111217
rect 252466 111143 252522 111152
rect 252284 111104 252336 111110
rect 252284 111046 252336 111052
rect 252098 108896 252154 108905
rect 252098 108831 252154 108840
rect 252192 107500 252244 107506
rect 252192 107442 252244 107448
rect 252204 105097 252232 107442
rect 252296 107001 252324 111046
rect 252376 110424 252428 110430
rect 252376 110366 252428 110372
rect 252388 109313 252416 110366
rect 252468 110356 252520 110362
rect 252468 110298 252520 110304
rect 252480 110265 252508 110298
rect 252466 110256 252522 110265
rect 252466 110191 252522 110200
rect 252374 109304 252430 109313
rect 252374 109239 252430 109248
rect 252376 108996 252428 109002
rect 252376 108938 252428 108944
rect 252388 107953 252416 108938
rect 252468 108928 252520 108934
rect 252468 108870 252520 108876
rect 252480 108361 252508 108870
rect 252466 108352 252522 108361
rect 252466 108287 252522 108296
rect 252374 107944 252430 107953
rect 252374 107879 252430 107888
rect 252376 107636 252428 107642
rect 252376 107578 252428 107584
rect 252282 106992 252338 107001
rect 252282 106927 252338 106936
rect 252388 106593 252416 107578
rect 252468 107568 252520 107574
rect 252466 107536 252468 107545
rect 252520 107536 252522 107545
rect 252466 107471 252522 107480
rect 252374 106584 252430 106593
rect 252374 106519 252430 106528
rect 252468 106276 252520 106282
rect 252468 106218 252520 106224
rect 252284 106208 252336 106214
rect 252284 106150 252336 106156
rect 252296 105641 252324 106150
rect 252480 106049 252508 106218
rect 252466 106040 252522 106049
rect 252466 105975 252522 105984
rect 252282 105632 252338 105641
rect 252282 105567 252338 105576
rect 252376 105596 252428 105602
rect 252376 105538 252428 105544
rect 252190 105088 252246 105097
rect 252190 105023 252246 105032
rect 252284 104780 252336 104786
rect 252284 104722 252336 104728
rect 252296 104145 252324 104722
rect 252282 104136 252338 104145
rect 252282 104071 252338 104080
rect 252006 103728 252062 103737
rect 252006 103663 252062 103672
rect 252192 102808 252244 102814
rect 252388 102785 252416 105538
rect 252468 104848 252520 104854
rect 252468 104790 252520 104796
rect 252480 104689 252508 104790
rect 252466 104680 252522 104689
rect 252466 104615 252522 104624
rect 252468 103488 252520 103494
rect 252468 103430 252520 103436
rect 252192 102750 252244 102756
rect 252374 102776 252430 102785
rect 251364 102128 251416 102134
rect 251364 102070 251416 102076
rect 251376 101833 251404 102070
rect 251362 101824 251418 101833
rect 251362 101759 251418 101768
rect 252204 100881 252232 102750
rect 252374 102711 252430 102720
rect 252480 102241 252508 103430
rect 252466 102232 252522 102241
rect 252466 102167 252522 102176
rect 252468 102060 252520 102066
rect 252468 102002 252520 102008
rect 252284 101448 252336 101454
rect 252480 101425 252508 102002
rect 252284 101390 252336 101396
rect 252466 101416 252522 101425
rect 252190 100872 252246 100881
rect 252190 100807 252246 100816
rect 252296 100473 252324 101390
rect 252466 101351 252522 101360
rect 252376 100700 252428 100706
rect 252376 100642 252428 100648
rect 252282 100464 252338 100473
rect 252282 100399 252338 100408
rect 252388 99521 252416 100642
rect 252468 100632 252520 100638
rect 252468 100574 252520 100580
rect 252480 99929 252508 100574
rect 252466 99920 252522 99929
rect 252466 99855 252522 99864
rect 252374 99512 252430 99521
rect 252374 99447 252430 99456
rect 252376 99340 252428 99346
rect 252376 99282 252428 99288
rect 251270 98560 251326 98569
rect 251270 98495 251326 98504
rect 252388 98025 252416 99282
rect 252468 99272 252520 99278
rect 252468 99214 252520 99220
rect 252480 98977 252508 99214
rect 252466 98968 252522 98977
rect 252466 98903 252522 98912
rect 252374 98016 252430 98025
rect 252374 97951 252430 97960
rect 252468 97980 252520 97986
rect 252468 97922 252520 97928
rect 252480 97617 252508 97922
rect 252466 97608 252522 97617
rect 252466 97543 252522 97552
rect 251270 97064 251326 97073
rect 251270 96999 251326 97008
rect 252466 97064 252522 97073
rect 252466 96999 252522 97008
rect 251178 96248 251234 96257
rect 251178 96183 251234 96192
rect 251192 93922 251220 96183
rect 251100 93894 251220 93922
rect 251100 93854 251128 93894
rect 251100 93826 251220 93854
rect 251192 91866 251220 93826
rect 251180 91860 251232 91866
rect 251180 91802 251232 91808
rect 251284 84194 251312 96999
rect 252480 96665 252508 96999
rect 252466 96656 252522 96665
rect 252466 96591 252522 96600
rect 251192 84166 251312 84194
rect 250444 11824 250496 11830
rect 250444 11766 250496 11772
rect 251192 9654 251220 84166
rect 253216 65618 253244 111794
rect 253308 102134 253336 143550
rect 253388 141432 253440 141438
rect 253388 141374 253440 141380
rect 253400 103358 253428 141374
rect 253480 137284 253532 137290
rect 253480 137226 253532 137232
rect 253492 125526 253520 137226
rect 253480 125520 253532 125526
rect 253480 125462 253532 125468
rect 254596 110294 254624 150418
rect 254676 146328 254728 146334
rect 254676 146270 254728 146276
rect 254584 110288 254636 110294
rect 254584 110230 254636 110236
rect 254688 107506 254716 146270
rect 255608 139398 255636 180202
rect 256700 176044 256752 176050
rect 256700 175986 256752 175992
rect 256712 170814 256740 175986
rect 256700 170808 256752 170814
rect 256700 170750 256752 170756
rect 256148 157616 256200 157622
rect 256148 157558 256200 157564
rect 256056 151836 256108 151842
rect 256056 151778 256108 151784
rect 255964 146396 256016 146402
rect 255964 146338 256016 146344
rect 255596 139392 255648 139398
rect 255596 139334 255648 139340
rect 254676 107500 254728 107506
rect 254676 107442 254728 107448
rect 255976 106214 256004 146338
rect 256068 111722 256096 151778
rect 256160 118590 256188 157558
rect 256804 150278 256832 183126
rect 256976 183116 257028 183122
rect 256976 183058 257028 183064
rect 256792 150272 256844 150278
rect 256792 150214 256844 150220
rect 256988 140690 257016 183058
rect 258092 169862 258120 199514
rect 259552 192500 259604 192506
rect 259552 192442 259604 192448
rect 259460 180396 259512 180402
rect 259460 180338 259512 180344
rect 258172 180328 258224 180334
rect 258172 180270 258224 180276
rect 258080 169856 258132 169862
rect 258080 169798 258132 169804
rect 258184 166258 258212 180270
rect 258264 178832 258316 178838
rect 258264 178774 258316 178780
rect 258276 167890 258304 178774
rect 258356 177404 258408 177410
rect 258356 177346 258408 177352
rect 258264 167884 258316 167890
rect 258264 167826 258316 167832
rect 258172 166252 258224 166258
rect 258172 166194 258224 166200
rect 258368 165782 258396 177346
rect 259472 171426 259500 180338
rect 259460 171420 259512 171426
rect 259460 171362 259512 171368
rect 259000 169788 259052 169794
rect 259000 169730 259052 169736
rect 258356 165776 258408 165782
rect 258356 165718 258408 165724
rect 258908 165640 258960 165646
rect 258908 165582 258960 165588
rect 258816 164280 258868 164286
rect 258816 164222 258868 164228
rect 258724 158772 258776 158778
rect 258724 158714 258776 158720
rect 257344 149728 257396 149734
rect 257344 149670 257396 149676
rect 256976 140684 257028 140690
rect 256976 140626 257028 140632
rect 256148 118584 256200 118590
rect 256148 118526 256200 118532
rect 256056 111716 256108 111722
rect 256056 111658 256108 111664
rect 255964 106208 256016 106214
rect 255964 106150 256016 106156
rect 253388 103352 253440 103358
rect 253388 103294 253440 103300
rect 253296 102128 253348 102134
rect 253296 102070 253348 102076
rect 257356 99278 257384 149670
rect 257436 140072 257488 140078
rect 257436 140014 257488 140020
rect 257448 104786 257476 140014
rect 258736 119474 258764 158714
rect 258828 126682 258856 164222
rect 258920 127498 258948 165582
rect 259012 142361 259040 169730
rect 259564 168978 259592 192442
rect 259644 188488 259696 188494
rect 259644 188430 259696 188436
rect 259656 172582 259684 188430
rect 259644 172576 259696 172582
rect 259644 172518 259696 172524
rect 259552 168972 259604 168978
rect 259552 168914 259604 168920
rect 259748 160818 259776 220118
rect 260932 211812 260984 211818
rect 260932 211754 260984 211760
rect 260840 178764 260892 178770
rect 260840 178706 260892 178712
rect 260288 171148 260340 171154
rect 260288 171090 260340 171096
rect 259736 160812 259788 160818
rect 259736 160754 259788 160760
rect 260104 160132 260156 160138
rect 260104 160074 260156 160080
rect 258998 142352 259054 142361
rect 258998 142287 259054 142296
rect 258908 127492 258960 127498
rect 258908 127434 258960 127440
rect 258816 126676 258868 126682
rect 258816 126618 258868 126624
rect 260116 120698 260144 160074
rect 260196 155984 260248 155990
rect 260196 155926 260248 155932
rect 260104 120692 260156 120698
rect 260104 120634 260156 120640
rect 258724 119468 258776 119474
rect 258724 119410 258776 119416
rect 260104 117360 260156 117366
rect 260104 117302 260156 117308
rect 257436 104780 257488 104786
rect 257436 104722 257488 104728
rect 257344 99272 257396 99278
rect 257344 99214 257396 99220
rect 258724 98048 258776 98054
rect 258724 97990 258776 97996
rect 255964 96688 256016 96694
rect 255964 96630 256016 96636
rect 253204 65612 253256 65618
rect 253204 65554 253256 65560
rect 255976 15910 256004 96630
rect 255964 15904 256016 15910
rect 255964 15846 256016 15852
rect 258736 14482 258764 97990
rect 258724 14476 258776 14482
rect 258724 14418 258776 14424
rect 251180 9648 251232 9654
rect 251180 9590 251232 9596
rect 177304 3528 177356 3534
rect 177304 3470 177356 3476
rect 235816 3528 235868 3534
rect 235816 3470 235868 3476
rect 238024 3528 238076 3534
rect 238024 3470 238076 3476
rect 235828 480 235856 3470
rect 260116 3466 260144 117302
rect 260208 116142 260236 155926
rect 260300 131578 260328 171090
rect 260852 169658 260880 178706
rect 260944 169726 260972 211754
rect 261116 203652 261168 203658
rect 261116 203594 261168 203600
rect 261024 180464 261076 180470
rect 261024 180406 261076 180412
rect 260932 169720 260984 169726
rect 260932 169662 260984 169668
rect 260840 169652 260892 169658
rect 260840 169594 260892 169600
rect 261036 168366 261064 180406
rect 261024 168360 261076 168366
rect 261024 168302 261076 168308
rect 261128 155854 261156 203594
rect 261576 168428 261628 168434
rect 261576 168370 261628 168376
rect 261484 162920 261536 162926
rect 261484 162862 261536 162868
rect 261116 155848 261168 155854
rect 261116 155790 261168 155796
rect 260288 131572 260340 131578
rect 260288 131514 260340 131520
rect 261496 124098 261524 162862
rect 261588 130422 261616 168370
rect 261668 167068 261720 167074
rect 261668 167010 261720 167016
rect 261576 130416 261628 130422
rect 261576 130358 261628 130364
rect 261680 129674 261708 167010
rect 262232 142118 262260 280230
rect 263600 247104 263652 247110
rect 263600 247046 263652 247052
rect 262312 198008 262364 198014
rect 262312 197950 262364 197956
rect 262324 146130 262352 197950
rect 262404 184340 262456 184346
rect 262404 184282 262456 184288
rect 262416 162722 262444 184282
rect 262496 182980 262548 182986
rect 262496 182922 262548 182928
rect 262508 165510 262536 182922
rect 263612 172378 263640 247046
rect 266372 238814 266400 697614
rect 283852 697610 283880 703520
rect 300136 700369 300164 703520
rect 305644 703112 305696 703118
rect 305644 703054 305696 703060
rect 300122 700360 300178 700369
rect 300122 700295 300178 700304
rect 283840 697604 283892 697610
rect 283840 697546 283892 697552
rect 286324 307828 286376 307834
rect 286324 307770 286376 307776
rect 267740 303680 267792 303686
rect 267740 303622 267792 303628
rect 266452 245676 266504 245682
rect 266452 245618 266504 245624
rect 266360 238808 266412 238814
rect 266360 238750 266412 238756
rect 264980 207800 265032 207806
rect 264980 207742 265032 207748
rect 263692 206372 263744 206378
rect 263692 206314 263744 206320
rect 263600 172372 263652 172378
rect 263600 172314 263652 172320
rect 262496 165504 262548 165510
rect 262496 165446 262548 165452
rect 263704 162790 263732 206314
rect 263784 177472 263836 177478
rect 263784 177414 263836 177420
rect 263692 162784 263744 162790
rect 263692 162726 263744 162732
rect 262404 162716 262456 162722
rect 262404 162658 262456 162664
rect 262956 158840 263008 158846
rect 262956 158782 263008 158788
rect 262864 156052 262916 156058
rect 262864 155994 262916 156000
rect 262312 146124 262364 146130
rect 262312 146066 262364 146072
rect 262220 142112 262272 142118
rect 262220 142054 262272 142060
rect 261668 129668 261720 129674
rect 261668 129610 261720 129616
rect 261484 124092 261536 124098
rect 261484 124034 261536 124040
rect 262876 117298 262904 155994
rect 262968 120018 262996 158782
rect 263796 157214 263824 177414
rect 264244 173936 264296 173942
rect 264244 173878 264296 173884
rect 263784 157208 263836 157214
rect 263784 157150 263836 157156
rect 264256 145586 264284 173878
rect 264992 165578 265020 207742
rect 266360 204944 266412 204950
rect 266360 204886 266412 204892
rect 265072 183048 265124 183054
rect 265072 182990 265124 182996
rect 264980 165572 265032 165578
rect 264980 165514 265032 165520
rect 265084 155922 265112 182990
rect 265808 171216 265860 171222
rect 265808 171158 265860 171164
rect 265716 169856 265768 169862
rect 265716 169798 265768 169804
rect 265072 155916 265124 155922
rect 265072 155858 265124 155864
rect 264520 154624 264572 154630
rect 264520 154566 264572 154572
rect 264336 150544 264388 150550
rect 264336 150486 264388 150492
rect 264244 145580 264296 145586
rect 264244 145522 264296 145528
rect 262956 120012 263008 120018
rect 262956 119954 263008 119960
rect 263048 119400 263100 119406
rect 263048 119342 263100 119348
rect 262864 117292 262916 117298
rect 262864 117234 262916 117240
rect 260196 116136 260248 116142
rect 260196 116078 260248 116084
rect 262864 109064 262916 109070
rect 262864 109006 262916 109012
rect 262876 26994 262904 109006
rect 263060 97986 263088 119342
rect 264244 114572 264296 114578
rect 264244 114514 264296 114520
rect 263048 97980 263100 97986
rect 263048 97922 263100 97928
rect 262864 26988 262916 26994
rect 262864 26930 262916 26936
rect 264256 25566 264284 114514
rect 264348 110362 264376 150486
rect 264428 147824 264480 147830
rect 264428 147766 264480 147772
rect 264336 110356 264388 110362
rect 264336 110298 264388 110304
rect 264440 107574 264468 147766
rect 264532 115938 264560 154566
rect 265622 145616 265678 145625
rect 265622 145551 265678 145560
rect 264520 115932 264572 115938
rect 264520 115874 264572 115880
rect 264428 107568 264480 107574
rect 264428 107510 264480 107516
rect 265636 104854 265664 145551
rect 265728 132394 265756 169798
rect 265820 138718 265848 171158
rect 266372 162858 266400 204886
rect 266360 162852 266412 162858
rect 266360 162794 266412 162800
rect 266464 144906 266492 245618
rect 267188 172576 267240 172582
rect 267188 172518 267240 172524
rect 267096 157480 267148 157486
rect 267096 157422 267148 157428
rect 266452 144900 266504 144906
rect 266452 144842 266504 144848
rect 265808 138712 265860 138718
rect 265808 138654 265860 138660
rect 267004 138100 267056 138106
rect 267004 138042 267056 138048
rect 265716 132388 265768 132394
rect 265716 132330 265768 132336
rect 265624 104848 265676 104854
rect 265624 104790 265676 104796
rect 264244 25560 264296 25566
rect 264244 25502 264296 25508
rect 267016 10402 267044 138042
rect 267108 118658 267136 157422
rect 267200 135182 267228 172518
rect 267752 164218 267780 303622
rect 281540 302320 281592 302326
rect 281540 302262 281592 302268
rect 280160 300892 280212 300898
rect 280160 300834 280212 300840
rect 277400 295452 277452 295458
rect 277400 295394 277452 295400
rect 270500 292664 270552 292670
rect 270500 292606 270552 292612
rect 267832 292596 267884 292602
rect 267832 292538 267884 292544
rect 267740 164212 267792 164218
rect 267740 164154 267792 164160
rect 267280 160744 267332 160750
rect 267280 160686 267332 160692
rect 267188 135176 267240 135182
rect 267188 135118 267240 135124
rect 267292 131034 267320 160686
rect 267844 160070 267872 292538
rect 269120 289876 269172 289882
rect 269120 289818 269172 289824
rect 267924 195356 267976 195362
rect 267924 195298 267976 195304
rect 267832 160064 267884 160070
rect 267832 160006 267884 160012
rect 267936 154494 267964 195298
rect 268384 174004 268436 174010
rect 268384 173946 268436 173952
rect 267924 154488 267976 154494
rect 267924 154430 267976 154436
rect 268396 136474 268424 173946
rect 268476 151904 268528 151910
rect 268476 151846 268528 151852
rect 268384 136468 268436 136474
rect 268384 136410 268436 136416
rect 267280 131028 267332 131034
rect 267280 130970 267332 130976
rect 268488 120766 268516 151846
rect 268568 143676 268620 143682
rect 268568 143618 268620 143624
rect 268476 120760 268528 120766
rect 268476 120702 268528 120708
rect 267096 118652 267148 118658
rect 267096 118594 267148 118600
rect 268384 117428 268436 117434
rect 268384 117370 268436 117376
rect 267188 116000 267240 116006
rect 267188 115942 267240 115948
rect 267096 103556 267148 103562
rect 267096 103498 267148 103504
rect 267108 39438 267136 103498
rect 267200 68338 267228 115942
rect 267188 68332 267240 68338
rect 267188 68274 267240 68280
rect 267096 39432 267148 39438
rect 267096 39374 267148 39380
rect 267004 10396 267056 10402
rect 267004 10338 267056 10344
rect 268396 4826 268424 117370
rect 268476 106480 268528 106486
rect 268476 106422 268528 106428
rect 268488 62830 268516 106422
rect 268580 103494 268608 143618
rect 269132 143478 269160 289818
rect 269212 189848 269264 189854
rect 269212 189790 269264 189796
rect 269224 153134 269252 189790
rect 269856 168496 269908 168502
rect 269856 168438 269908 168444
rect 269764 162988 269816 162994
rect 269764 162930 269816 162936
rect 269212 153128 269264 153134
rect 269212 153070 269264 153076
rect 269120 143472 269172 143478
rect 269120 143414 269172 143420
rect 269776 124166 269804 162930
rect 269868 129742 269896 168438
rect 270512 143546 270540 292606
rect 276664 266484 276716 266490
rect 276664 266426 276716 266432
rect 273260 254040 273312 254046
rect 273260 253982 273312 253988
rect 271880 210520 271932 210526
rect 271880 210462 271932 210468
rect 270684 209092 270736 209098
rect 270684 209034 270736 209040
rect 270592 188420 270644 188426
rect 270592 188362 270644 188368
rect 270500 143540 270552 143546
rect 270500 143482 270552 143488
rect 269948 142180 270000 142186
rect 269948 142122 270000 142128
rect 269856 129736 269908 129742
rect 269856 129678 269908 129684
rect 269764 124160 269816 124166
rect 269764 124102 269816 124108
rect 269764 120148 269816 120154
rect 269764 120090 269816 120096
rect 268568 103488 268620 103494
rect 268568 103430 268620 103436
rect 268476 62824 268528 62830
rect 268476 62766 268528 62772
rect 269776 43518 269804 120090
rect 269960 102814 269988 142122
rect 270604 136542 270632 188362
rect 270696 157282 270724 209034
rect 271328 167136 271380 167142
rect 271328 167078 271380 167084
rect 270684 157276 270736 157282
rect 270684 157218 270736 157224
rect 270592 136536 270644 136542
rect 270592 136478 270644 136484
rect 271144 131164 271196 131170
rect 271144 131106 271196 131112
rect 269948 102808 270000 102814
rect 269948 102750 270000 102756
rect 269856 102196 269908 102202
rect 269856 102138 269908 102144
rect 269764 43512 269816 43518
rect 269764 43454 269816 43460
rect 269868 35290 269896 102138
rect 271156 49026 271184 131106
rect 271340 128246 271368 167078
rect 271892 137834 271920 210462
rect 271972 200796 272024 200802
rect 271972 200738 272024 200744
rect 271984 154562 272012 200738
rect 272616 165708 272668 165714
rect 272616 165650 272668 165656
rect 271972 154556 272024 154562
rect 271972 154498 272024 154504
rect 271880 137828 271932 137834
rect 271880 137770 271932 137776
rect 271328 128240 271380 128246
rect 271328 128182 271380 128188
rect 272524 127084 272576 127090
rect 272524 127026 272576 127032
rect 271236 127016 271288 127022
rect 271236 126958 271288 126964
rect 271248 53106 271276 126958
rect 272536 75206 272564 127026
rect 272628 126954 272656 165650
rect 273272 150346 273300 253982
rect 276020 231192 276072 231198
rect 276020 231134 276072 231140
rect 273352 216028 273404 216034
rect 273352 215970 273404 215976
rect 273260 150340 273312 150346
rect 273260 150282 273312 150288
rect 273364 146266 273392 215970
rect 273444 194064 273496 194070
rect 273444 194006 273496 194012
rect 273352 146260 273404 146266
rect 273352 146202 273404 146208
rect 273456 146198 273484 194006
rect 274732 188624 274784 188630
rect 274732 188566 274784 188572
rect 274640 187060 274692 187066
rect 274640 187002 274692 187008
rect 274088 164348 274140 164354
rect 274088 164290 274140 164296
rect 273444 146192 273496 146198
rect 273444 146134 273496 146140
rect 273996 129804 274048 129810
rect 273996 129746 274048 129752
rect 272616 126948 272668 126954
rect 272616 126890 272668 126896
rect 273904 125656 273956 125662
rect 273904 125598 273956 125604
rect 272524 75200 272576 75206
rect 272524 75142 272576 75148
rect 271236 53100 271288 53106
rect 271236 53042 271288 53048
rect 271144 49020 271196 49026
rect 271144 48962 271196 48968
rect 273916 44878 273944 125598
rect 274008 55962 274036 129746
rect 274100 125594 274128 164290
rect 274652 140758 274680 187002
rect 274744 147626 274772 188566
rect 276032 151774 276060 231134
rect 276112 199504 276164 199510
rect 276112 199446 276164 199452
rect 276020 151768 276072 151774
rect 276020 151710 276072 151716
rect 276124 148986 276152 199446
rect 276676 182986 276704 266426
rect 276664 182980 276716 182986
rect 276664 182922 276716 182928
rect 276664 172644 276716 172650
rect 276664 172586 276716 172592
rect 276112 148980 276164 148986
rect 276112 148922 276164 148928
rect 274732 147620 274784 147626
rect 274732 147562 274784 147568
rect 275284 140956 275336 140962
rect 275284 140898 275336 140904
rect 274640 140752 274692 140758
rect 274640 140694 274692 140700
rect 274088 125588 274140 125594
rect 274088 125530 274140 125536
rect 275296 104174 275324 140898
rect 276676 135250 276704 172586
rect 277412 137902 277440 295394
rect 278780 209160 278832 209166
rect 278780 209102 278832 209108
rect 277492 207732 277544 207738
rect 277492 207674 277544 207680
rect 277504 137970 277532 207674
rect 278792 150414 278820 209102
rect 278780 150408 278832 150414
rect 278780 150350 278832 150356
rect 280172 149054 280200 300834
rect 280804 165776 280856 165782
rect 280804 165718 280856 165724
rect 280160 149048 280212 149054
rect 280160 148990 280212 148996
rect 280816 142866 280844 165718
rect 281552 157350 281580 302262
rect 284944 267776 284996 267782
rect 284944 267718 284996 267724
rect 284956 177342 284984 267718
rect 284944 177336 284996 177342
rect 286336 177313 286364 307770
rect 302884 306400 302936 306406
rect 302884 306342 302936 306348
rect 287704 305040 287756 305046
rect 287704 304982 287756 304988
rect 287716 179382 287744 304982
rect 289084 244384 289136 244390
rect 289084 244326 289136 244332
rect 289096 184346 289124 244326
rect 298744 217388 298796 217394
rect 298744 217330 298796 217336
rect 289084 184340 289136 184346
rect 289084 184282 289136 184288
rect 287704 179376 287756 179382
rect 287704 179318 287756 179324
rect 298756 178809 298784 217330
rect 300124 215960 300176 215966
rect 300124 215902 300176 215908
rect 300136 181626 300164 215902
rect 300124 181620 300176 181626
rect 300124 181562 300176 181568
rect 302896 178945 302924 306342
rect 305656 238746 305684 703054
rect 332520 702545 332548 703520
rect 348804 703050 348832 703520
rect 348792 703044 348844 703050
rect 348792 702986 348844 702992
rect 332506 702536 332562 702545
rect 332506 702471 332562 702480
rect 364996 699718 365024 703520
rect 397472 702846 397500 703520
rect 413664 702982 413692 703520
rect 413652 702976 413704 702982
rect 413652 702918 413704 702924
rect 397460 702840 397512 702846
rect 397460 702782 397512 702788
rect 429856 702710 429884 703520
rect 462332 702914 462360 703520
rect 462320 702908 462372 702914
rect 462320 702850 462372 702856
rect 478524 702778 478552 703520
rect 494808 703118 494836 703520
rect 494796 703112 494848 703118
rect 494796 703054 494848 703060
rect 478512 702772 478564 702778
rect 478512 702714 478564 702720
rect 429844 702704 429896 702710
rect 429844 702646 429896 702652
rect 527192 702642 527220 703520
rect 527180 702636 527232 702642
rect 527180 702578 527232 702584
rect 543476 702434 543504 703520
rect 559668 702574 559696 703520
rect 559656 702568 559708 702574
rect 559656 702510 559708 702516
rect 580908 702500 580960 702506
rect 580908 702442 580960 702448
rect 542372 702406 543504 702434
rect 359464 699712 359516 699718
rect 359464 699654 359516 699660
rect 364984 699712 365036 699718
rect 364984 699654 365036 699660
rect 334624 302252 334676 302258
rect 334624 302194 334676 302200
rect 325792 299600 325844 299606
rect 325792 299542 325844 299548
rect 308404 296948 308456 296954
rect 308404 296890 308456 296896
rect 307024 294092 307076 294098
rect 307024 294034 307076 294040
rect 305644 238740 305696 238746
rect 305644 238682 305696 238688
rect 305644 225616 305696 225622
rect 305644 225558 305696 225564
rect 304264 220108 304316 220114
rect 304264 220050 304316 220056
rect 302882 178936 302938 178945
rect 302882 178871 302938 178880
rect 298742 178800 298798 178809
rect 298742 178735 298798 178744
rect 304276 177410 304304 220050
rect 304264 177404 304316 177410
rect 304264 177346 304316 177352
rect 284944 177278 284996 177284
rect 286322 177304 286378 177313
rect 286322 177239 286378 177248
rect 305656 176662 305684 225558
rect 307036 181490 307064 294034
rect 307024 181484 307076 181490
rect 307024 181426 307076 181432
rect 305644 176656 305696 176662
rect 305644 176598 305696 176604
rect 307114 175264 307170 175273
rect 307114 175199 307170 175208
rect 306562 174856 306618 174865
rect 306562 174791 306618 174800
rect 287796 174072 287848 174078
rect 287796 174014 287848 174020
rect 284944 172712 284996 172718
rect 284944 172654 284996 172660
rect 282276 167204 282328 167210
rect 282276 167146 282328 167152
rect 281540 157344 281592 157350
rect 281540 157286 281592 157292
rect 281080 149116 281132 149122
rect 281080 149058 281132 149064
rect 280804 142860 280856 142866
rect 280804 142802 280856 142808
rect 280988 142248 281040 142254
rect 280988 142190 281040 142196
rect 279516 139460 279568 139466
rect 279516 139402 279568 139408
rect 277492 137964 277544 137970
rect 277492 137906 277544 137912
rect 277400 137896 277452 137902
rect 277400 137838 277452 137844
rect 278136 135312 278188 135318
rect 278136 135254 278188 135260
rect 276664 135244 276716 135250
rect 276664 135186 276716 135192
rect 276756 133952 276808 133958
rect 276756 133894 276808 133900
rect 276664 128376 276716 128382
rect 276664 128318 276716 128324
rect 275376 124976 275428 124982
rect 275376 124918 275428 124924
rect 275388 108934 275416 124918
rect 275376 108928 275428 108934
rect 275376 108870 275428 108876
rect 275284 104168 275336 104174
rect 275284 104110 275336 104116
rect 275284 102264 275336 102270
rect 275284 102206 275336 102212
rect 273996 55956 274048 55962
rect 273996 55898 274048 55904
rect 273904 44872 273956 44878
rect 273904 44814 273956 44820
rect 269856 35284 269908 35290
rect 269856 35226 269908 35232
rect 275296 7614 275324 102206
rect 276676 17270 276704 128318
rect 276768 50386 276796 133894
rect 278044 131232 278096 131238
rect 278044 131174 278096 131180
rect 276756 50380 276808 50386
rect 276756 50322 276808 50328
rect 278056 22778 278084 131174
rect 278148 47598 278176 135254
rect 279424 103624 279476 103630
rect 279424 103566 279476 103572
rect 278136 47592 278188 47598
rect 278136 47534 278188 47540
rect 278044 22772 278096 22778
rect 278044 22714 278096 22720
rect 276664 17264 276716 17270
rect 276664 17206 276716 17212
rect 279436 13122 279464 103566
rect 279528 76634 279556 139402
rect 280804 138168 280856 138174
rect 280804 138110 280856 138116
rect 279516 76628 279568 76634
rect 279516 76570 279568 76576
rect 279424 13116 279476 13122
rect 279424 13058 279476 13064
rect 275284 7608 275336 7614
rect 275284 7550 275336 7556
rect 268384 4820 268436 4826
rect 268384 4762 268436 4768
rect 260104 3460 260156 3466
rect 260104 3402 260156 3408
rect 280816 2174 280844 138110
rect 280896 116068 280948 116074
rect 280896 116010 280948 116016
rect 280908 24138 280936 116010
rect 281000 102066 281028 142190
rect 281092 116618 281120 149058
rect 282184 132524 282236 132530
rect 282184 132466 282236 132472
rect 281080 116612 281132 116618
rect 281080 116554 281132 116560
rect 280988 102060 281040 102066
rect 280988 102002 281040 102008
rect 280896 24132 280948 24138
rect 280896 24074 280948 24080
rect 282196 8974 282224 132466
rect 282288 128314 282316 167146
rect 282460 153264 282512 153270
rect 282460 153206 282512 153212
rect 282276 128308 282328 128314
rect 282276 128250 282328 128256
rect 282368 122868 282420 122874
rect 282368 122810 282420 122816
rect 282276 107908 282328 107914
rect 282276 107850 282328 107856
rect 282288 18630 282316 107850
rect 282380 61402 282408 122810
rect 282472 115258 282500 153206
rect 283564 135380 283616 135386
rect 283564 135322 283616 135328
rect 282460 115252 282512 115258
rect 282460 115194 282512 115200
rect 282368 61396 282420 61402
rect 282368 61338 282420 61344
rect 283576 38010 283604 135322
rect 284956 133822 284984 172654
rect 286416 169924 286468 169930
rect 286416 169866 286468 169872
rect 286324 161560 286376 161566
rect 286324 161502 286376 161508
rect 285036 154692 285088 154698
rect 285036 154634 285088 154640
rect 284944 133816 284996 133822
rect 284944 133758 284996 133764
rect 285048 114442 285076 154634
rect 285220 145580 285272 145586
rect 285220 145522 285272 145528
rect 285128 129872 285180 129878
rect 285128 129814 285180 129820
rect 285036 114436 285088 114442
rect 285036 114378 285088 114384
rect 284944 113212 284996 113218
rect 284944 113154 284996 113160
rect 283656 100768 283708 100774
rect 283656 100710 283708 100716
rect 283564 38004 283616 38010
rect 283564 37946 283616 37952
rect 283668 28286 283696 100710
rect 283656 28280 283708 28286
rect 283656 28222 283708 28228
rect 282276 18624 282328 18630
rect 282276 18566 282328 18572
rect 282184 8968 282236 8974
rect 282184 8910 282236 8916
rect 284956 6186 284984 113154
rect 285036 104916 285088 104922
rect 285036 104858 285088 104864
rect 285048 14550 285076 104858
rect 285140 40730 285168 129814
rect 285232 106282 285260 145522
rect 286336 122738 286364 161502
rect 286428 132462 286456 169866
rect 287808 136610 287836 174014
rect 306576 173942 306604 174791
rect 306564 173936 306616 173942
rect 306564 173878 306616 173884
rect 306562 172272 306618 172281
rect 306562 172207 306618 172216
rect 306576 171290 306604 172207
rect 289176 171284 289228 171290
rect 289176 171226 289228 171232
rect 306564 171284 306616 171290
rect 306564 171226 306616 171232
rect 287980 150612 288032 150618
rect 287980 150554 288032 150560
rect 287796 136604 287848 136610
rect 287796 136546 287848 136552
rect 287704 135448 287756 135454
rect 287704 135390 287756 135396
rect 286600 133204 286652 133210
rect 286600 133146 286652 133152
rect 286416 132456 286468 132462
rect 286416 132398 286468 132404
rect 286508 125724 286560 125730
rect 286508 125666 286560 125672
rect 286324 122732 286376 122738
rect 286324 122674 286376 122680
rect 286416 121508 286468 121514
rect 286416 121450 286468 121456
rect 285220 106276 285272 106282
rect 285220 106218 285272 106224
rect 286324 98116 286376 98122
rect 286324 98058 286376 98064
rect 285128 40724 285180 40730
rect 285128 40666 285180 40672
rect 285036 14544 285088 14550
rect 285036 14486 285088 14492
rect 286336 11762 286364 98058
rect 286428 44946 286456 121450
rect 286520 69698 286548 125666
rect 286612 99346 286640 133146
rect 286600 99340 286652 99346
rect 286600 99282 286652 99288
rect 286508 69692 286560 69698
rect 286508 69634 286560 69640
rect 286416 44940 286468 44946
rect 286416 44882 286468 44888
rect 287716 43450 287744 135390
rect 287888 114640 287940 114646
rect 287888 114582 287940 114588
rect 287796 109132 287848 109138
rect 287796 109074 287848 109080
rect 287704 43444 287756 43450
rect 287704 43386 287756 43392
rect 287808 22846 287836 109074
rect 287900 65550 287928 114582
rect 287992 110430 288020 150554
rect 289084 139528 289136 139534
rect 289084 139470 289136 139476
rect 287980 110424 288032 110430
rect 287980 110366 288032 110372
rect 287888 65544 287940 65550
rect 287888 65486 287940 65492
rect 287796 22840 287848 22846
rect 287796 22782 287848 22788
rect 286324 11756 286376 11762
rect 286324 11698 286376 11704
rect 289096 10334 289124 139470
rect 289188 133890 289216 171226
rect 306562 170640 306618 170649
rect 306562 170575 306618 170584
rect 306576 169930 306604 170575
rect 306564 169924 306616 169930
rect 306564 169866 306616 169872
rect 291844 168564 291896 168570
rect 291844 168506 291896 168512
rect 289360 161628 289412 161634
rect 289360 161570 289412 161576
rect 289176 133884 289228 133890
rect 289176 133826 289228 133832
rect 289176 127152 289228 127158
rect 289176 127094 289228 127100
rect 289188 51746 289216 127094
rect 289372 122670 289400 161570
rect 290648 146940 290700 146946
rect 290648 146882 290700 146888
rect 290556 132592 290608 132598
rect 290556 132534 290608 132540
rect 289360 122664 289412 122670
rect 289360 122606 289412 122612
rect 289268 121576 289320 121582
rect 289268 121518 289320 121524
rect 289280 53174 289308 121518
rect 290464 120216 290516 120222
rect 290464 120158 290516 120164
rect 289360 96756 289412 96762
rect 289360 96698 289412 96704
rect 289268 53168 289320 53174
rect 289268 53110 289320 53116
rect 289176 51740 289228 51746
rect 289176 51682 289228 51688
rect 289372 31074 289400 96698
rect 290476 42158 290504 120158
rect 290568 58750 290596 132534
rect 290660 121446 290688 146882
rect 291856 131102 291884 168506
rect 307022 165064 307078 165073
rect 307022 164999 307078 165008
rect 300400 164416 300452 164422
rect 300400 164358 300452 164364
rect 297456 163056 297508 163062
rect 297456 162998 297508 163004
rect 295984 157548 296036 157554
rect 295984 157490 296036 157496
rect 292120 145648 292172 145654
rect 292120 145590 292172 145596
rect 291936 134020 291988 134026
rect 291936 133962 291988 133968
rect 291844 131096 291896 131102
rect 291844 131038 291896 131044
rect 290648 121440 290700 121446
rect 290648 121382 290700 121388
rect 291844 120284 291896 120290
rect 291844 120226 291896 120232
rect 290648 99408 290700 99414
rect 290648 99350 290700 99356
rect 290556 58744 290608 58750
rect 290556 58686 290608 58692
rect 290464 42152 290516 42158
rect 290464 42094 290516 42100
rect 290660 36582 290688 99350
rect 291856 40798 291884 120226
rect 291948 57254 291976 133962
rect 292028 122936 292080 122942
rect 292028 122878 292080 122884
rect 291936 57248 291988 57254
rect 291936 57190 291988 57196
rect 292040 50454 292068 122878
rect 292132 109002 292160 145590
rect 294880 140888 294932 140894
rect 294880 140830 294932 140836
rect 293224 136672 293276 136678
rect 293224 136614 293276 136620
rect 292120 108996 292172 109002
rect 292120 108938 292172 108944
rect 292212 107772 292264 107778
rect 292212 107714 292264 107720
rect 292224 76566 292252 107714
rect 292212 76560 292264 76566
rect 292212 76502 292264 76508
rect 292028 50448 292080 50454
rect 292028 50390 292080 50396
rect 291844 40792 291896 40798
rect 291844 40734 291896 40740
rect 290648 36576 290700 36582
rect 290648 36518 290700 36524
rect 293236 33862 293264 136614
rect 294788 131300 294840 131306
rect 294788 131242 294840 131248
rect 293316 117496 293368 117502
rect 293316 117438 293368 117444
rect 293328 35222 293356 117438
rect 293408 114708 293460 114714
rect 293408 114650 293460 114656
rect 293420 66910 293448 114650
rect 294604 113280 294656 113286
rect 294604 113222 294656 113228
rect 293408 66904 293460 66910
rect 293408 66846 293460 66852
rect 293316 35216 293368 35222
rect 293316 35158 293368 35164
rect 293224 33856 293276 33862
rect 293224 33798 293276 33804
rect 289360 31068 289412 31074
rect 289360 31010 289412 31016
rect 294616 19990 294644 113222
rect 294696 102332 294748 102338
rect 294696 102274 294748 102280
rect 294708 29646 294736 102274
rect 294800 73846 294828 131242
rect 294892 100638 294920 140830
rect 295996 137358 296024 157490
rect 296168 156120 296220 156126
rect 296168 156062 296220 156068
rect 295984 137352 296036 137358
rect 295984 137294 296036 137300
rect 296076 128444 296128 128450
rect 296076 128386 296128 128392
rect 295984 124228 296036 124234
rect 295984 124170 296036 124176
rect 294880 100632 294932 100638
rect 294880 100574 294932 100580
rect 294788 73840 294840 73846
rect 294788 73782 294840 73788
rect 294696 29640 294748 29646
rect 294696 29582 294748 29588
rect 294604 19984 294656 19990
rect 294604 19926 294656 19932
rect 289084 10328 289136 10334
rect 289084 10270 289136 10276
rect 284944 6180 284996 6186
rect 284944 6122 284996 6128
rect 280804 2168 280856 2174
rect 280804 2110 280856 2116
rect 295996 2106 296024 124170
rect 296088 21418 296116 128386
rect 296180 117978 296208 156062
rect 297364 136740 297416 136746
rect 297364 136682 297416 136688
rect 296260 129940 296312 129946
rect 296260 129882 296312 129888
rect 296168 117972 296220 117978
rect 296168 117914 296220 117920
rect 296168 116136 296220 116142
rect 296168 116078 296220 116084
rect 296180 33794 296208 116078
rect 296272 71058 296300 129882
rect 296260 71052 296312 71058
rect 296260 70994 296312 71000
rect 296168 33788 296220 33794
rect 296168 33730 296220 33736
rect 296076 21412 296128 21418
rect 296076 21354 296128 21360
rect 297376 7682 297404 136682
rect 297468 124914 297496 162998
rect 298744 158908 298796 158914
rect 298744 158850 298796 158856
rect 297456 124908 297508 124914
rect 297456 124850 297508 124856
rect 297548 121644 297600 121650
rect 297548 121586 297600 121592
rect 297456 99476 297508 99482
rect 297456 99418 297508 99424
rect 297468 26926 297496 99418
rect 297560 51814 297588 121586
rect 298756 120086 298784 158850
rect 300216 154760 300268 154766
rect 300216 154702 300268 154708
rect 299112 149796 299164 149802
rect 299112 149738 299164 149744
rect 299020 143744 299072 143750
rect 299020 143686 299072 143692
rect 298928 124296 298980 124302
rect 298928 124238 298980 124244
rect 298744 120080 298796 120086
rect 298744 120022 298796 120028
rect 298836 118856 298888 118862
rect 298836 118798 298888 118804
rect 298744 104984 298796 104990
rect 298744 104926 298796 104932
rect 297548 51808 297600 51814
rect 297548 51750 297600 51756
rect 297456 26920 297508 26926
rect 297456 26862 297508 26868
rect 298756 15978 298784 104926
rect 298848 39370 298876 118798
rect 298940 72554 298968 124238
rect 299032 105602 299060 143686
rect 299124 113150 299152 149738
rect 300124 125792 300176 125798
rect 300124 125734 300176 125740
rect 299112 113144 299164 113150
rect 299112 113086 299164 113092
rect 299020 105596 299072 105602
rect 299020 105538 299072 105544
rect 299020 100836 299072 100842
rect 299020 100778 299072 100784
rect 298928 72548 298980 72554
rect 298928 72490 298980 72496
rect 299032 58682 299060 100778
rect 299020 58676 299072 58682
rect 299020 58618 299072 58624
rect 300136 46238 300164 125734
rect 300228 114510 300256 154702
rect 300308 142316 300360 142322
rect 300308 142258 300360 142264
rect 300216 114504 300268 114510
rect 300216 114446 300268 114452
rect 300216 110560 300268 110566
rect 300216 110502 300268 110508
rect 300228 66978 300256 110502
rect 300320 101454 300348 142258
rect 300412 126274 300440 164358
rect 304540 160200 304592 160206
rect 304540 160142 304592 160148
rect 303528 153332 303580 153338
rect 303528 153274 303580 153280
rect 303540 148345 303568 153274
rect 304264 151972 304316 151978
rect 304264 151914 304316 151920
rect 303526 148336 303582 148345
rect 303526 148271 303582 148280
rect 301780 147688 301832 147694
rect 301780 147630 301832 147636
rect 301596 128512 301648 128518
rect 301596 128454 301648 128460
rect 300400 126268 300452 126274
rect 300400 126210 300452 126216
rect 301504 111920 301556 111926
rect 301504 111862 301556 111868
rect 300492 105052 300544 105058
rect 300492 104994 300544 105000
rect 300308 101448 300360 101454
rect 300308 101390 300360 101396
rect 300400 100904 300452 100910
rect 300400 100846 300452 100852
rect 300216 66972 300268 66978
rect 300216 66914 300268 66920
rect 300412 64190 300440 100846
rect 300504 72486 300532 104994
rect 300492 72480 300544 72486
rect 300492 72422 300544 72428
rect 300400 64184 300452 64190
rect 300400 64126 300452 64132
rect 300124 46232 300176 46238
rect 300124 46174 300176 46180
rect 298836 39364 298888 39370
rect 298836 39306 298888 39312
rect 301516 25634 301544 111862
rect 301608 42090 301636 128454
rect 301688 118720 301740 118726
rect 301688 118662 301740 118668
rect 301700 55894 301728 118662
rect 301792 111110 301820 147630
rect 302884 135516 302936 135522
rect 302884 135458 302936 135464
rect 301780 111104 301832 111110
rect 301780 111046 301832 111052
rect 301688 55888 301740 55894
rect 301688 55830 301740 55836
rect 301596 42084 301648 42090
rect 301596 42026 301648 42032
rect 302896 36650 302924 135458
rect 303068 124364 303120 124370
rect 303068 124306 303120 124312
rect 302976 107704 303028 107710
rect 302976 107646 303028 107652
rect 302884 36644 302936 36650
rect 302884 36586 302936 36592
rect 301504 25628 301556 25634
rect 301504 25570 301556 25576
rect 302988 21486 303016 107646
rect 303080 75274 303108 124306
rect 304276 111790 304304 151914
rect 304448 140820 304500 140826
rect 304448 140762 304500 140768
rect 304356 123004 304408 123010
rect 304356 122946 304408 122952
rect 304264 111784 304316 111790
rect 304264 111726 304316 111732
rect 303160 110492 303212 110498
rect 303160 110434 303212 110440
rect 303068 75268 303120 75274
rect 303068 75210 303120 75216
rect 303172 68406 303200 110434
rect 304264 106412 304316 106418
rect 304264 106354 304316 106360
rect 303160 68400 303212 68406
rect 303160 68342 303212 68348
rect 302976 21480 303028 21486
rect 302976 21422 303028 21428
rect 304276 17338 304304 106354
rect 304368 49094 304396 122946
rect 304460 100706 304488 140762
rect 304552 123486 304580 160142
rect 306562 159080 306618 159089
rect 306562 159015 306618 159024
rect 306576 158914 306604 159015
rect 306564 158908 306616 158914
rect 306564 158850 306616 158856
rect 306930 158264 306986 158273
rect 306930 158199 306986 158208
rect 306944 157622 306972 158199
rect 306932 157616 306984 157622
rect 306932 157558 306984 157564
rect 305734 157448 305790 157457
rect 305734 157383 305790 157392
rect 305642 145072 305698 145081
rect 305642 145007 305698 145016
rect 304540 123480 304592 123486
rect 304540 123422 304592 123428
rect 305656 112470 305684 145007
rect 305748 129062 305776 157383
rect 306562 154864 306618 154873
rect 306562 154799 306618 154808
rect 306576 154698 306604 154799
rect 306564 154692 306616 154698
rect 306564 154634 306616 154640
rect 306562 154456 306618 154465
rect 306562 154391 306618 154400
rect 306576 153270 306604 154391
rect 306564 153264 306616 153270
rect 306564 153206 306616 153212
rect 306654 153232 306710 153241
rect 306654 153167 306710 153176
rect 306668 149802 306696 153167
rect 306930 151056 306986 151065
rect 306930 150991 306986 151000
rect 306944 150482 306972 150991
rect 306932 150476 306984 150482
rect 306932 150418 306984 150424
rect 306656 149796 306708 149802
rect 306656 149738 306708 149744
rect 306562 148880 306618 148889
rect 306562 148815 306618 148824
rect 305918 147928 305974 147937
rect 305918 147863 305974 147872
rect 305736 129056 305788 129062
rect 305736 128998 305788 129004
rect 305826 118824 305882 118833
rect 305826 118759 305882 118768
rect 305644 112464 305696 112470
rect 305644 112406 305696 112412
rect 305642 110664 305698 110673
rect 305642 110599 305698 110608
rect 304540 109200 304592 109206
rect 304540 109142 304592 109148
rect 304448 100700 304500 100706
rect 304448 100642 304500 100648
rect 304552 71126 304580 109142
rect 304540 71120 304592 71126
rect 304540 71062 304592 71068
rect 304356 49088 304408 49094
rect 304356 49030 304408 49036
rect 305656 24206 305684 110599
rect 305734 106720 305790 106729
rect 305734 106655 305790 106664
rect 305748 28354 305776 106655
rect 305840 64258 305868 118759
rect 305932 107642 305960 147863
rect 306576 147830 306604 148815
rect 306564 147824 306616 147830
rect 306564 147766 306616 147772
rect 306930 146840 306986 146849
rect 306930 146775 306986 146784
rect 306944 146334 306972 146775
rect 306932 146328 306984 146334
rect 306932 146270 306984 146276
rect 306562 143440 306618 143449
rect 306562 143375 306618 143384
rect 306576 142254 306604 143375
rect 306564 142248 306616 142254
rect 306564 142190 306616 142196
rect 306562 142080 306618 142089
rect 306562 142015 306618 142024
rect 306576 140894 306604 142015
rect 306564 140888 306616 140894
rect 306564 140830 306616 140836
rect 306746 140856 306802 140865
rect 306746 140791 306802 140800
rect 306562 139088 306618 139097
rect 306562 139023 306618 139032
rect 306576 138038 306604 139023
rect 306564 138032 306616 138038
rect 306564 137974 306616 137980
rect 306562 136232 306618 136241
rect 306562 136167 306618 136176
rect 306576 135454 306604 136167
rect 306564 135448 306616 135454
rect 306564 135390 306616 135396
rect 306760 133210 306788 140791
rect 306930 140040 306986 140049
rect 306930 139975 306986 139984
rect 306944 139534 306972 139975
rect 306932 139528 306984 139534
rect 306932 139470 306984 139476
rect 307036 137290 307064 164999
rect 307128 149734 307156 175199
rect 307574 174448 307630 174457
rect 307574 174383 307630 174392
rect 307588 174078 307616 174383
rect 307576 174072 307628 174078
rect 307576 174014 307628 174020
rect 307666 174040 307722 174049
rect 307666 173975 307668 173984
rect 307720 173975 307722 173984
rect 307668 173946 307720 173952
rect 307574 173632 307630 173641
rect 307574 173567 307630 173576
rect 307484 172712 307536 172718
rect 307482 172680 307484 172689
rect 307536 172680 307538 172689
rect 307588 172650 307616 173567
rect 307666 173224 307722 173233
rect 307666 173159 307722 173168
rect 307482 172615 307538 172624
rect 307576 172644 307628 172650
rect 307576 172586 307628 172592
rect 307680 172582 307708 173159
rect 307668 172576 307720 172582
rect 307668 172518 307720 172524
rect 307574 171864 307630 171873
rect 307574 171799 307630 171808
rect 307588 171222 307616 171799
rect 307666 171456 307722 171465
rect 307666 171391 307722 171400
rect 307576 171216 307628 171222
rect 307576 171158 307628 171164
rect 307680 171154 307708 171391
rect 307668 171148 307720 171154
rect 307668 171090 307720 171096
rect 307574 171048 307630 171057
rect 307574 170983 307630 170992
rect 307588 169862 307616 170983
rect 307666 170232 307722 170241
rect 307666 170167 307722 170176
rect 307576 169856 307628 169862
rect 307390 169824 307446 169833
rect 307576 169798 307628 169804
rect 307680 169794 307708 170167
rect 307390 169759 307446 169768
rect 307668 169788 307720 169794
rect 307298 166424 307354 166433
rect 307298 166359 307354 166368
rect 307312 165714 307340 166359
rect 307300 165708 307352 165714
rect 307300 165650 307352 165656
rect 307298 165472 307354 165481
rect 307298 165407 307354 165416
rect 307312 164286 307340 165407
rect 307300 164280 307352 164286
rect 307300 164222 307352 164228
rect 307404 161474 307432 169759
rect 307668 169730 307720 169736
rect 307666 169280 307722 169289
rect 307666 169215 307722 169224
rect 307574 168872 307630 168881
rect 307574 168807 307630 168816
rect 307484 168496 307536 168502
rect 307482 168464 307484 168473
rect 307536 168464 307538 168473
rect 307588 168434 307616 168807
rect 307680 168570 307708 169215
rect 307668 168564 307720 168570
rect 307668 168506 307720 168512
rect 307482 168399 307538 168408
rect 307576 168428 307628 168434
rect 307576 168370 307628 168376
rect 307482 168056 307538 168065
rect 307482 167991 307538 168000
rect 307496 167074 307524 167991
rect 307574 167648 307630 167657
rect 307574 167583 307630 167592
rect 307588 167142 307616 167583
rect 307666 167240 307722 167249
rect 307666 167175 307668 167184
rect 307720 167175 307722 167184
rect 307668 167146 307720 167152
rect 307576 167136 307628 167142
rect 307576 167078 307628 167084
rect 307484 167068 307536 167074
rect 307484 167010 307536 167016
rect 307574 166832 307630 166841
rect 307574 166767 307630 166776
rect 307588 165646 307616 166767
rect 307666 165880 307722 165889
rect 307666 165815 307722 165824
rect 307680 165782 307708 165815
rect 307668 165776 307720 165782
rect 307668 165718 307720 165724
rect 307576 165640 307628 165646
rect 307576 165582 307628 165588
rect 307666 164656 307722 164665
rect 307666 164591 307722 164600
rect 307576 164416 307628 164422
rect 307576 164358 307628 164364
rect 307588 164257 307616 164358
rect 307680 164354 307708 164591
rect 307668 164348 307720 164354
rect 307668 164290 307720 164296
rect 307574 164248 307630 164257
rect 307574 164183 307630 164192
rect 307574 163840 307630 163849
rect 307574 163775 307630 163784
rect 307482 163432 307538 163441
rect 307482 163367 307538 163376
rect 307496 162994 307524 163367
rect 307588 163062 307616 163775
rect 307576 163056 307628 163062
rect 307576 162998 307628 163004
rect 307666 163024 307722 163033
rect 307484 162988 307536 162994
rect 307666 162959 307722 162968
rect 307484 162930 307536 162936
rect 307680 162926 307708 162959
rect 307668 162920 307720 162926
rect 307668 162862 307720 162868
rect 307574 162480 307630 162489
rect 307574 162415 307630 162424
rect 307482 162072 307538 162081
rect 307482 162007 307538 162016
rect 307496 161498 307524 162007
rect 307588 161634 307616 162415
rect 307666 161664 307722 161673
rect 307576 161628 307628 161634
rect 307666 161599 307722 161608
rect 307576 161570 307628 161576
rect 307680 161566 307708 161599
rect 307668 161560 307720 161566
rect 307668 161502 307720 161508
rect 307312 161446 307432 161474
rect 307484 161492 307536 161498
rect 307206 160848 307262 160857
rect 307206 160783 307262 160792
rect 307116 149728 307168 149734
rect 307116 149670 307168 149676
rect 307220 146946 307248 160783
rect 307312 160750 307340 161446
rect 307484 161434 307536 161440
rect 307574 161256 307630 161265
rect 307574 161191 307630 161200
rect 307300 160744 307352 160750
rect 307300 160686 307352 160692
rect 307588 160138 307616 161191
rect 307666 160440 307722 160449
rect 307666 160375 307722 160384
rect 307680 160206 307708 160375
rect 307668 160200 307720 160206
rect 307668 160142 307720 160148
rect 307576 160132 307628 160138
rect 307576 160074 307628 160080
rect 307298 160032 307354 160041
rect 307298 159967 307354 159976
rect 307312 158846 307340 159967
rect 307666 159624 307722 159633
rect 307666 159559 307722 159568
rect 307300 158840 307352 158846
rect 307300 158782 307352 158788
rect 307680 158778 307708 159559
rect 307668 158772 307720 158778
rect 307668 158714 307720 158720
rect 307574 158672 307630 158681
rect 307574 158607 307630 158616
rect 307588 157486 307616 158607
rect 307666 157856 307722 157865
rect 307666 157791 307722 157800
rect 307680 157554 307708 157791
rect 307668 157548 307720 157554
rect 307668 157490 307720 157496
rect 307576 157480 307628 157486
rect 307576 157422 307628 157428
rect 307482 157040 307538 157049
rect 307482 156975 307538 156984
rect 307496 156058 307524 156975
rect 307574 156632 307630 156641
rect 307574 156567 307630 156576
rect 307484 156052 307536 156058
rect 307484 155994 307536 156000
rect 307588 155990 307616 156567
rect 307666 156224 307722 156233
rect 307666 156159 307722 156168
rect 307680 156126 307708 156159
rect 307668 156120 307720 156126
rect 307668 156062 307720 156068
rect 307576 155984 307628 155990
rect 307576 155926 307628 155932
rect 307298 155680 307354 155689
rect 307298 155615 307354 155624
rect 307312 154630 307340 155615
rect 307666 155272 307722 155281
rect 307666 155207 307722 155216
rect 307680 154766 307708 155207
rect 307668 154760 307720 154766
rect 307668 154702 307720 154708
rect 307300 154624 307352 154630
rect 307300 154566 307352 154572
rect 307666 153640 307722 153649
rect 307666 153575 307722 153584
rect 307680 153338 307708 153575
rect 307668 153332 307720 153338
rect 307668 153274 307720 153280
rect 307482 152688 307538 152697
rect 307482 152623 307538 152632
rect 307496 151842 307524 152623
rect 307574 152280 307630 152289
rect 307574 152215 307630 152224
rect 307588 151978 307616 152215
rect 307576 151972 307628 151978
rect 307576 151914 307628 151920
rect 307668 151904 307720 151910
rect 307666 151872 307668 151881
rect 307720 151872 307722 151881
rect 307484 151836 307536 151842
rect 307666 151807 307722 151816
rect 307484 151778 307536 151784
rect 307298 151464 307354 151473
rect 307298 151399 307354 151408
rect 307312 150550 307340 151399
rect 307666 150648 307722 150657
rect 307666 150583 307668 150592
rect 307720 150583 307722 150592
rect 307668 150554 307720 150560
rect 307300 150544 307352 150550
rect 307300 150486 307352 150492
rect 307666 150240 307722 150249
rect 307666 150175 307722 150184
rect 307390 149832 307446 149841
rect 307390 149767 307446 149776
rect 307298 147248 307354 147257
rect 307298 147183 307354 147192
rect 307208 146940 307260 146946
rect 307208 146882 307260 146888
rect 307312 146402 307340 147183
rect 307300 146396 307352 146402
rect 307300 146338 307352 146344
rect 307114 145888 307170 145897
rect 307114 145823 307170 145832
rect 307128 140078 307156 145823
rect 307404 145014 307432 149767
rect 307574 149288 307630 149297
rect 307574 149223 307630 149232
rect 307482 147656 307538 147665
rect 307482 147591 307538 147600
rect 307496 145586 307524 147591
rect 307588 145654 307616 149223
rect 307680 149122 307708 150175
rect 307668 149116 307720 149122
rect 307668 149058 307720 149064
rect 307666 148472 307722 148481
rect 307666 148407 307722 148416
rect 307680 147694 307708 148407
rect 307668 147688 307720 147694
rect 307668 147630 307720 147636
rect 307576 145648 307628 145654
rect 307576 145590 307628 145596
rect 307484 145580 307536 145586
rect 307484 145522 307536 145528
rect 307312 144986 307432 145014
rect 307312 142154 307340 144986
rect 307390 144936 307446 144945
rect 307390 144871 307446 144880
rect 307404 143562 307432 144871
rect 307482 144664 307538 144673
rect 307482 144599 307538 144608
rect 307496 143750 307524 144599
rect 307574 144256 307630 144265
rect 307574 144191 307630 144200
rect 307484 143744 307536 143750
rect 307484 143686 307536 143692
rect 307588 143682 307616 144191
rect 307666 143848 307722 143857
rect 307666 143783 307722 143792
rect 307576 143676 307628 143682
rect 307576 143618 307628 143624
rect 307680 143614 307708 143783
rect 307668 143608 307720 143614
rect 307404 143534 307524 143562
rect 307668 143550 307720 143556
rect 307312 142126 307432 142154
rect 307206 140448 307262 140457
rect 307206 140383 307262 140392
rect 307116 140072 307168 140078
rect 307116 140014 307168 140020
rect 307114 137864 307170 137873
rect 307114 137799 307170 137808
rect 307024 137284 307076 137290
rect 307024 137226 307076 137232
rect 306748 133204 306800 133210
rect 306748 133146 306800 133152
rect 306746 128888 306802 128897
rect 306746 128823 306802 128832
rect 306760 128518 306788 128823
rect 306748 128512 306800 128518
rect 306748 128454 306800 128460
rect 306930 125080 306986 125089
rect 306930 125015 306986 125024
rect 306944 124370 306972 125015
rect 306932 124364 306984 124370
rect 306932 124306 306984 124312
rect 306562 118688 306618 118697
rect 306562 118623 306618 118632
rect 306576 117366 306604 118623
rect 306564 117360 306616 117366
rect 306564 117302 306616 117308
rect 306746 116648 306802 116657
rect 306746 116583 306802 116592
rect 306760 116006 306788 116583
rect 306748 116000 306800 116006
rect 306748 115942 306800 115948
rect 306010 107672 306066 107681
rect 305920 107636 305972 107642
rect 306010 107607 306066 107616
rect 305920 107578 305972 107584
rect 306024 73914 306052 107607
rect 306930 103048 306986 103057
rect 306930 102983 306986 102992
rect 306944 102338 306972 102983
rect 306932 102332 306984 102338
rect 306932 102274 306984 102280
rect 307022 98696 307078 98705
rect 307022 98631 307078 98640
rect 306932 96756 306984 96762
rect 306932 96698 306984 96704
rect 306944 96665 306972 96698
rect 306930 96656 306986 96665
rect 306930 96591 306986 96600
rect 306012 73908 306064 73914
rect 306012 73850 306064 73856
rect 305828 64252 305880 64258
rect 305828 64194 305880 64200
rect 307036 37942 307064 98631
rect 307128 89010 307156 137799
rect 307220 135250 307248 140383
rect 307298 139632 307354 139641
rect 307298 139567 307354 139576
rect 307312 139466 307340 139567
rect 307300 139460 307352 139466
rect 307300 139402 307352 139408
rect 307298 135688 307354 135697
rect 307298 135623 307354 135632
rect 307312 135522 307340 135623
rect 307300 135516 307352 135522
rect 307300 135458 307352 135464
rect 307208 135244 307260 135250
rect 307208 135186 307260 135192
rect 307206 132696 307262 132705
rect 307206 132631 307262 132640
rect 307220 90370 307248 132631
rect 307404 132494 307432 142126
rect 307496 141438 307524 143534
rect 307574 143032 307630 143041
rect 307574 142967 307630 142976
rect 307588 142186 307616 142967
rect 307666 142488 307722 142497
rect 307666 142423 307722 142432
rect 307680 142322 307708 142423
rect 307668 142316 307720 142322
rect 307668 142258 307720 142264
rect 307576 142180 307628 142186
rect 307576 142122 307628 142128
rect 307574 141672 307630 141681
rect 307574 141607 307630 141616
rect 307484 141432 307536 141438
rect 307484 141374 307536 141380
rect 307588 140826 307616 141607
rect 307666 141264 307722 141273
rect 307666 141199 307722 141208
rect 307680 140962 307708 141199
rect 307668 140956 307720 140962
rect 307668 140898 307720 140904
rect 307576 140820 307628 140826
rect 307576 140762 307628 140768
rect 307574 138680 307630 138689
rect 307574 138615 307630 138624
rect 307588 138106 307616 138615
rect 307666 138272 307722 138281
rect 307666 138207 307722 138216
rect 307680 138174 307708 138207
rect 307668 138168 307720 138174
rect 307668 138110 307720 138116
rect 307576 138100 307628 138106
rect 307576 138042 307628 138048
rect 307574 137456 307630 137465
rect 307574 137391 307630 137400
rect 307588 136678 307616 137391
rect 307666 137048 307722 137057
rect 307666 136983 307722 136992
rect 307680 136746 307708 136983
rect 307668 136740 307720 136746
rect 307668 136682 307720 136688
rect 307576 136672 307628 136678
rect 307482 136640 307538 136649
rect 307576 136614 307628 136620
rect 307482 136575 307538 136584
rect 307496 135386 307524 136575
rect 307484 135380 307536 135386
rect 307484 135322 307536 135328
rect 307668 135312 307720 135318
rect 307666 135280 307668 135289
rect 307720 135280 307722 135289
rect 307484 135244 307536 135250
rect 307666 135215 307722 135224
rect 307484 135186 307536 135192
rect 307312 132466 307432 132494
rect 307312 124982 307340 132466
rect 307390 132288 307446 132297
rect 307390 132223 307446 132232
rect 307404 131238 307432 132223
rect 307392 131232 307444 131238
rect 307392 131174 307444 131180
rect 307496 129962 307524 135186
rect 307574 134872 307630 134881
rect 307574 134807 307630 134816
rect 307588 134026 307616 134807
rect 307666 134464 307722 134473
rect 307666 134399 307722 134408
rect 307576 134020 307628 134026
rect 307576 133962 307628 133968
rect 307680 133958 307708 134399
rect 307668 133952 307720 133958
rect 307668 133894 307720 133900
rect 307574 133648 307630 133657
rect 307574 133583 307630 133592
rect 307588 132530 307616 133583
rect 307666 133240 307722 133249
rect 307666 133175 307722 133184
rect 307680 132598 307708 133175
rect 307668 132592 307720 132598
rect 307668 132534 307720 132540
rect 307576 132524 307628 132530
rect 307576 132466 307628 132472
rect 307574 131880 307630 131889
rect 307574 131815 307630 131824
rect 307588 131170 307616 131815
rect 307666 131472 307722 131481
rect 307666 131407 307722 131416
rect 307680 131306 307708 131407
rect 307668 131300 307720 131306
rect 307668 131242 307720 131248
rect 307576 131164 307628 131170
rect 307576 131106 307628 131112
rect 307666 131064 307722 131073
rect 307666 130999 307722 131008
rect 307404 129934 307524 129962
rect 307574 129976 307630 129985
rect 307300 124976 307352 124982
rect 307300 124918 307352 124924
rect 307298 124672 307354 124681
rect 307298 124607 307354 124616
rect 307312 91798 307340 124607
rect 307404 119406 307432 129934
rect 307680 129946 307708 130999
rect 307574 129911 307630 129920
rect 307668 129940 307720 129946
rect 307484 129872 307536 129878
rect 307482 129840 307484 129849
rect 307536 129840 307538 129849
rect 307588 129810 307616 129911
rect 307668 129882 307720 129888
rect 307482 129775 307538 129784
rect 307576 129804 307628 129810
rect 307576 129746 307628 129752
rect 307574 129296 307630 129305
rect 307574 129231 307630 129240
rect 307588 128382 307616 129231
rect 307666 128480 307722 128489
rect 307666 128415 307668 128424
rect 307720 128415 307722 128424
rect 307668 128386 307720 128392
rect 307576 128376 307628 128382
rect 307576 128318 307628 128324
rect 307482 128072 307538 128081
rect 307482 128007 307538 128016
rect 307496 127022 307524 128007
rect 307574 127664 307630 127673
rect 307574 127599 307630 127608
rect 307588 127090 307616 127599
rect 307666 127256 307722 127265
rect 307666 127191 307722 127200
rect 307680 127158 307708 127191
rect 307668 127152 307720 127158
rect 307668 127094 307720 127100
rect 307576 127084 307628 127090
rect 307576 127026 307628 127032
rect 307484 127016 307536 127022
rect 307484 126958 307536 126964
rect 307482 126848 307538 126857
rect 307482 126783 307538 126792
rect 307496 125662 307524 126783
rect 307574 126440 307630 126449
rect 307574 126375 307630 126384
rect 307588 125730 307616 126375
rect 307666 125896 307722 125905
rect 307666 125831 307722 125840
rect 307680 125798 307708 125831
rect 307668 125792 307720 125798
rect 307668 125734 307720 125740
rect 307576 125724 307628 125730
rect 307576 125666 307628 125672
rect 307484 125656 307536 125662
rect 307484 125598 307536 125604
rect 307574 125488 307630 125497
rect 307574 125423 307630 125432
rect 307588 124302 307616 125423
rect 307576 124296 307628 124302
rect 307576 124238 307628 124244
rect 307666 124264 307722 124273
rect 307666 124199 307668 124208
rect 307720 124199 307722 124208
rect 307668 124170 307720 124176
rect 307482 123856 307538 123865
rect 307482 123791 307538 123800
rect 307496 122942 307524 123791
rect 307666 123448 307722 123457
rect 307666 123383 307722 123392
rect 307574 123040 307630 123049
rect 307680 123010 307708 123383
rect 307574 122975 307630 122984
rect 307668 123004 307720 123010
rect 307484 122936 307536 122942
rect 307484 122878 307536 122884
rect 307588 122874 307616 122975
rect 307668 122946 307720 122952
rect 307576 122868 307628 122874
rect 307576 122810 307628 122816
rect 307482 122496 307538 122505
rect 307482 122431 307538 122440
rect 307496 121514 307524 122431
rect 307574 122088 307630 122097
rect 307574 122023 307630 122032
rect 307588 121650 307616 122023
rect 307666 121680 307722 121689
rect 307576 121644 307628 121650
rect 307666 121615 307722 121624
rect 307576 121586 307628 121592
rect 307680 121582 307708 121615
rect 307668 121576 307720 121582
rect 307668 121518 307720 121524
rect 307484 121508 307536 121514
rect 307484 121450 307536 121456
rect 307482 121272 307538 121281
rect 307482 121207 307538 121216
rect 307496 120154 307524 121207
rect 307574 120864 307630 120873
rect 307574 120799 307630 120808
rect 307588 120222 307616 120799
rect 307666 120456 307722 120465
rect 307666 120391 307722 120400
rect 307680 120290 307708 120391
rect 307668 120284 307720 120290
rect 307668 120226 307720 120232
rect 307576 120216 307628 120222
rect 307576 120158 307628 120164
rect 307484 120148 307536 120154
rect 307484 120090 307536 120096
rect 307482 120048 307538 120057
rect 307482 119983 307538 119992
rect 307392 119400 307444 119406
rect 307392 119342 307444 119348
rect 307496 118726 307524 119983
rect 307574 119640 307630 119649
rect 307574 119575 307630 119584
rect 307588 118833 307616 119575
rect 307666 119096 307722 119105
rect 307666 119031 307722 119040
rect 307680 118862 307708 119031
rect 307668 118856 307720 118862
rect 307574 118824 307630 118833
rect 307668 118798 307720 118804
rect 307574 118759 307630 118768
rect 307484 118720 307536 118726
rect 307484 118662 307536 118668
rect 307574 117872 307630 117881
rect 307574 117807 307630 117816
rect 307588 117434 307616 117807
rect 307668 117496 307720 117502
rect 307666 117464 307668 117473
rect 307720 117464 307722 117473
rect 307576 117428 307628 117434
rect 307666 117399 307722 117408
rect 307576 117370 307628 117376
rect 307574 117056 307630 117065
rect 307574 116991 307630 117000
rect 307588 116142 307616 116991
rect 307666 116240 307722 116249
rect 307666 116175 307722 116184
rect 307576 116136 307628 116142
rect 307576 116078 307628 116084
rect 307680 116074 307708 116175
rect 307668 116068 307720 116074
rect 307668 116010 307720 116016
rect 307482 115696 307538 115705
rect 307482 115631 307538 115640
rect 307496 114578 307524 115631
rect 307574 115288 307630 115297
rect 307574 115223 307630 115232
rect 307588 114714 307616 115223
rect 307666 114880 307722 114889
rect 307666 114815 307722 114824
rect 307576 114708 307628 114714
rect 307576 114650 307628 114656
rect 307680 114646 307708 114815
rect 307668 114640 307720 114646
rect 307668 114582 307720 114588
rect 307484 114572 307536 114578
rect 307484 114514 307536 114520
rect 307666 113656 307722 113665
rect 307666 113591 307722 113600
rect 307680 113286 307708 113591
rect 307668 113280 307720 113286
rect 307574 113248 307630 113257
rect 307668 113222 307720 113228
rect 307574 113183 307576 113192
rect 307628 113183 307630 113192
rect 307576 113154 307628 113160
rect 307666 112024 307722 112033
rect 307666 111959 307722 111968
rect 307484 111920 307536 111926
rect 307482 111888 307484 111897
rect 307536 111888 307538 111897
rect 307680 111858 307708 111959
rect 307482 111823 307538 111832
rect 307668 111852 307720 111858
rect 307668 111794 307720 111800
rect 307574 111480 307630 111489
rect 307574 111415 307630 111424
rect 307588 110566 307616 111415
rect 307666 111072 307722 111081
rect 307666 111007 307722 111016
rect 307576 110560 307628 110566
rect 307576 110502 307628 110508
rect 307680 110498 307708 111007
rect 307668 110492 307720 110498
rect 307668 110434 307720 110440
rect 307482 110256 307538 110265
rect 307482 110191 307538 110200
rect 307496 109206 307524 110191
rect 307574 109848 307630 109857
rect 307574 109783 307630 109792
rect 307484 109200 307536 109206
rect 307484 109142 307536 109148
rect 307588 109138 307616 109783
rect 307666 109304 307722 109313
rect 307666 109239 307722 109248
rect 307576 109132 307628 109138
rect 307576 109074 307628 109080
rect 307680 109070 307708 109239
rect 307668 109064 307720 109070
rect 307668 109006 307720 109012
rect 307482 108896 307538 108905
rect 307482 108831 307538 108840
rect 307496 107681 307524 108831
rect 307666 108488 307722 108497
rect 307666 108423 307722 108432
rect 307574 108080 307630 108089
rect 307574 108015 307630 108024
rect 307588 107710 307616 108015
rect 307680 107914 307708 108423
rect 307668 107908 307720 107914
rect 307668 107850 307720 107856
rect 307668 107772 307720 107778
rect 307668 107714 307720 107720
rect 307576 107704 307628 107710
rect 307482 107672 307538 107681
rect 307680 107681 307708 107714
rect 307576 107646 307628 107652
rect 307666 107672 307722 107681
rect 307482 107607 307538 107616
rect 307666 107607 307722 107616
rect 307666 107264 307722 107273
rect 307666 107199 307722 107208
rect 307484 106480 307536 106486
rect 307482 106448 307484 106457
rect 307536 106448 307538 106457
rect 307680 106418 307708 107199
rect 307482 106383 307538 106392
rect 307668 106412 307720 106418
rect 307668 106354 307720 106360
rect 307482 105904 307538 105913
rect 307482 105839 307538 105848
rect 307496 104990 307524 105839
rect 307666 105496 307722 105505
rect 307666 105431 307722 105440
rect 307574 105088 307630 105097
rect 307680 105058 307708 105431
rect 307574 105023 307630 105032
rect 307668 105052 307720 105058
rect 307484 104984 307536 104990
rect 307484 104926 307536 104932
rect 307588 104922 307616 105023
rect 307668 104994 307720 105000
rect 307576 104916 307628 104922
rect 307576 104858 307628 104864
rect 307574 104680 307630 104689
rect 307574 104615 307630 104624
rect 307588 103562 307616 104615
rect 307666 103864 307722 103873
rect 307666 103799 307722 103808
rect 307680 103630 307708 103799
rect 307668 103624 307720 103630
rect 307668 103566 307720 103572
rect 307576 103556 307628 103562
rect 307576 103498 307628 103504
rect 307574 103456 307630 103465
rect 307574 103391 307630 103400
rect 307588 102270 307616 103391
rect 307666 102504 307722 102513
rect 307666 102439 307722 102448
rect 307576 102264 307628 102270
rect 307576 102206 307628 102212
rect 307680 102202 307708 102439
rect 307668 102196 307720 102202
rect 307668 102138 307720 102144
rect 307482 101688 307538 101697
rect 307482 101623 307538 101632
rect 307496 100842 307524 101623
rect 307574 101280 307630 101289
rect 307574 101215 307630 101224
rect 307588 100910 307616 101215
rect 307576 100904 307628 100910
rect 307576 100846 307628 100852
rect 307666 100872 307722 100881
rect 307484 100836 307536 100842
rect 307666 100807 307722 100816
rect 307484 100778 307536 100784
rect 307680 100774 307708 100807
rect 307668 100768 307720 100774
rect 307668 100710 307720 100716
rect 307574 100464 307630 100473
rect 307574 100399 307630 100408
rect 307588 99482 307616 100399
rect 307666 100056 307722 100065
rect 307666 99991 307722 100000
rect 307576 99476 307628 99482
rect 307576 99418 307628 99424
rect 307680 99414 307708 99991
rect 307668 99408 307720 99414
rect 307668 99350 307720 99356
rect 307574 99104 307630 99113
rect 307574 99039 307630 99048
rect 307588 98122 307616 99039
rect 307666 98288 307722 98297
rect 307666 98223 307722 98232
rect 307576 98116 307628 98122
rect 307576 98058 307628 98064
rect 307680 98054 307708 98223
rect 307668 98048 307720 98054
rect 307668 97990 307720 97996
rect 307666 97472 307722 97481
rect 307666 97407 307722 97416
rect 307680 96694 307708 97407
rect 307668 96688 307720 96694
rect 307668 96630 307720 96636
rect 307666 96248 307722 96257
rect 307666 96183 307722 96192
rect 307680 95266 307708 96183
rect 307668 95260 307720 95266
rect 307668 95202 307720 95208
rect 308416 95130 308444 296890
rect 322938 292632 322994 292641
rect 322938 292567 322994 292576
rect 321560 280220 321612 280226
rect 321560 280162 321612 280168
rect 313924 278792 313976 278798
rect 313924 278734 313976 278740
rect 309784 265056 309836 265062
rect 309784 264998 309836 265004
rect 308496 184272 308548 184278
rect 308496 184214 308548 184220
rect 308508 96626 308536 184214
rect 309138 114472 309194 114481
rect 309138 114407 309194 114416
rect 309152 113121 309180 114407
rect 309138 113112 309194 113121
rect 309138 113047 309194 113056
rect 308496 96620 308548 96626
rect 308496 96562 308548 96568
rect 308404 95124 308456 95130
rect 308404 95066 308456 95072
rect 309796 95062 309824 264998
rect 312544 239420 312596 239426
rect 312544 239362 312596 239368
rect 312556 177546 312584 239362
rect 312544 177540 312596 177546
rect 312544 177482 312596 177488
rect 313936 175982 313964 278734
rect 316684 252612 316736 252618
rect 316684 252554 316736 252560
rect 315304 228472 315356 228478
rect 315304 228414 315356 228420
rect 315316 177478 315344 228414
rect 316696 181694 316724 252554
rect 318064 242276 318116 242282
rect 318064 242218 318116 242224
rect 316684 181688 316736 181694
rect 316684 181630 316736 181636
rect 318076 181558 318104 242218
rect 320824 235340 320876 235346
rect 320824 235282 320876 235288
rect 320836 190454 320864 235282
rect 320836 190426 321324 190454
rect 316316 181552 316368 181558
rect 316316 181494 316368 181500
rect 318064 181552 318116 181558
rect 318064 181494 318116 181500
rect 315304 177472 315356 177478
rect 315304 177414 315356 177420
rect 316038 176760 316094 176769
rect 316038 176695 316094 176704
rect 313924 175976 313976 175982
rect 316052 175930 316080 176695
rect 316328 176225 316356 181494
rect 316314 176216 316370 176225
rect 316314 176151 316370 176160
rect 313924 175918 313976 175924
rect 316020 175902 316080 175930
rect 321296 169697 321324 190426
rect 321468 176656 321520 176662
rect 321468 176598 321520 176604
rect 321480 176089 321508 176598
rect 321466 176080 321522 176089
rect 321466 176015 321522 176024
rect 321468 175976 321520 175982
rect 321468 175918 321520 175924
rect 321480 175273 321508 175918
rect 321466 175264 321522 175273
rect 321466 175199 321522 175208
rect 321282 169688 321338 169697
rect 321282 169623 321338 169632
rect 321572 124273 321600 280162
rect 321652 217320 321704 217326
rect 321652 217262 321704 217268
rect 321664 127537 321692 217262
rect 321744 191344 321796 191350
rect 321744 191286 321796 191292
rect 321756 148345 321784 191286
rect 322952 157049 322980 292567
rect 325698 290592 325754 290601
rect 325698 290527 325754 290536
rect 324596 261520 324648 261526
rect 324596 261462 324648 261468
rect 323124 214600 323176 214606
rect 323124 214542 323176 214548
rect 323032 199436 323084 199442
rect 323032 199378 323084 199384
rect 322938 157040 322994 157049
rect 322938 156975 322994 156984
rect 321742 148336 321798 148345
rect 321742 148271 321798 148280
rect 321650 127528 321706 127537
rect 321650 127463 321706 127472
rect 321558 124264 321614 124273
rect 321558 124199 321614 124208
rect 321558 105088 321614 105097
rect 321558 105023 321614 105032
rect 321282 98832 321338 98841
rect 321282 98767 321338 98776
rect 321296 95169 321324 98767
rect 321374 97336 321430 97345
rect 321374 97271 321430 97280
rect 321282 95160 321338 95169
rect 321282 95095 321338 95104
rect 321388 95062 321416 97271
rect 321466 96656 321522 96665
rect 321466 96591 321468 96600
rect 321520 96591 321522 96600
rect 321468 96562 321520 96568
rect 309784 95056 309836 95062
rect 309784 94998 309836 95004
rect 321376 95056 321428 95062
rect 321376 94998 321428 95004
rect 321572 93702 321600 105023
rect 321650 103728 321706 103737
rect 321650 103663 321706 103672
rect 321664 93838 321692 103663
rect 323044 103193 323072 199378
rect 323136 121689 323164 214542
rect 324412 193996 324464 194002
rect 324412 193938 324464 193944
rect 323216 184204 323268 184210
rect 323216 184146 323268 184152
rect 323228 165481 323256 184146
rect 324320 172508 324372 172514
rect 324320 172450 324372 172456
rect 324332 172417 324360 172450
rect 324318 172408 324374 172417
rect 324318 172343 324374 172352
rect 324320 171080 324372 171086
rect 324320 171022 324372 171028
rect 324332 170921 324360 171022
rect 324318 170912 324374 170921
rect 324318 170847 324374 170856
rect 324424 168609 324452 193938
rect 324504 185768 324556 185774
rect 324504 185710 324556 185716
rect 324516 174049 324544 185710
rect 324502 174040 324558 174049
rect 324502 173975 324558 173984
rect 324608 173233 324636 261462
rect 324594 173224 324650 173233
rect 324594 173159 324650 173168
rect 324410 168600 324466 168609
rect 324410 168535 324466 168544
rect 324320 168360 324372 168366
rect 324320 168302 324372 168308
rect 324332 167793 324360 168302
rect 324412 168292 324464 168298
rect 324412 168234 324464 168240
rect 324318 167784 324374 167793
rect 324318 167719 324374 167728
rect 324424 167113 324452 168234
rect 324410 167104 324466 167113
rect 324410 167039 324466 167048
rect 324320 167000 324372 167006
rect 324320 166942 324372 166948
rect 324332 166297 324360 166942
rect 324318 166288 324374 166297
rect 324318 166223 324374 166232
rect 324320 165572 324372 165578
rect 324320 165514 324372 165520
rect 323214 165472 323270 165481
rect 323214 165407 323270 165416
rect 324332 164801 324360 165514
rect 324318 164792 324374 164801
rect 324318 164727 324374 164736
rect 324412 164212 324464 164218
rect 324412 164154 324464 164160
rect 324320 164144 324372 164150
rect 324320 164086 324372 164092
rect 324332 163985 324360 164086
rect 324318 163976 324374 163985
rect 324318 163911 324374 163920
rect 324424 163169 324452 164154
rect 324410 163160 324466 163169
rect 324410 163095 324466 163104
rect 324320 162852 324372 162858
rect 324320 162794 324372 162800
rect 324332 162489 324360 162794
rect 324318 162480 324374 162489
rect 324318 162415 324374 162424
rect 324320 161900 324372 161906
rect 324320 161842 324372 161848
rect 324332 161673 324360 161842
rect 324318 161664 324374 161673
rect 324318 161599 324374 161608
rect 324320 161424 324372 161430
rect 324320 161366 324372 161372
rect 324332 160857 324360 161366
rect 324412 161356 324464 161362
rect 324412 161298 324464 161304
rect 324318 160848 324374 160857
rect 324318 160783 324374 160792
rect 324424 160177 324452 161298
rect 324410 160168 324466 160177
rect 324410 160103 324466 160112
rect 324320 160064 324372 160070
rect 324320 160006 324372 160012
rect 324332 159361 324360 160006
rect 324318 159352 324374 159361
rect 324318 159287 324374 159296
rect 324412 158704 324464 158710
rect 324412 158646 324464 158652
rect 324320 158636 324372 158642
rect 324320 158578 324372 158584
rect 324332 158545 324360 158578
rect 324318 158536 324374 158545
rect 324318 158471 324374 158480
rect 324424 157865 324452 158646
rect 324410 157856 324466 157865
rect 324410 157791 324466 157800
rect 324320 157344 324372 157350
rect 324320 157286 324372 157292
rect 324332 156369 324360 157286
rect 324318 156360 324374 156369
rect 324318 156295 324374 156304
rect 324412 155916 324464 155922
rect 324412 155858 324464 155864
rect 324320 155848 324372 155854
rect 324320 155790 324372 155796
rect 324332 155553 324360 155790
rect 324318 155544 324374 155553
rect 324318 155479 324374 155488
rect 324424 154737 324452 155858
rect 324410 154728 324466 154737
rect 324410 154663 324466 154672
rect 324320 154556 324372 154562
rect 324320 154498 324372 154504
rect 324332 154057 324360 154498
rect 324318 154048 324374 154057
rect 324318 153983 324374 153992
rect 324320 153808 324372 153814
rect 324320 153750 324372 153756
rect 324332 153241 324360 153750
rect 324318 153232 324374 153241
rect 324318 153167 324374 153176
rect 324412 153196 324464 153202
rect 324412 153138 324464 153144
rect 324424 152425 324452 153138
rect 324410 152416 324466 152425
rect 324410 152351 324466 152360
rect 324318 151736 324374 151745
rect 324318 151671 324320 151680
rect 324372 151671 324374 151680
rect 324320 151642 324372 151648
rect 324320 150408 324372 150414
rect 324320 150350 324372 150356
rect 324332 150113 324360 150350
rect 324412 150272 324464 150278
rect 324412 150214 324464 150220
rect 324318 150104 324374 150113
rect 324318 150039 324374 150048
rect 324424 149433 324452 150214
rect 324410 149424 324466 149433
rect 324410 149359 324466 149368
rect 324320 149048 324372 149054
rect 324320 148990 324372 148996
rect 324332 148617 324360 148990
rect 324318 148608 324374 148617
rect 324318 148543 324374 148552
rect 324320 147620 324372 147626
rect 324320 147562 324372 147568
rect 324332 147121 324360 147562
rect 324318 147112 324374 147121
rect 324318 147047 324374 147056
rect 324318 146296 324374 146305
rect 324318 146231 324320 146240
rect 324372 146231 324374 146240
rect 324320 146202 324372 146208
rect 324412 146192 324464 146198
rect 324412 146134 324464 146140
rect 324424 145489 324452 146134
rect 324410 145480 324466 145489
rect 324410 145415 324466 145424
rect 324320 144900 324372 144906
rect 324320 144842 324372 144848
rect 324332 144809 324360 144842
rect 324412 144832 324464 144838
rect 324318 144800 324374 144809
rect 324412 144774 324464 144780
rect 324318 144735 324374 144744
rect 324424 143993 324452 144774
rect 324410 143984 324466 143993
rect 324410 143919 324466 143928
rect 324412 143540 324464 143546
rect 324412 143482 324464 143488
rect 324320 143472 324372 143478
rect 324320 143414 324372 143420
rect 324332 143177 324360 143414
rect 324318 143168 324374 143177
rect 324318 143103 324374 143112
rect 324424 142497 324452 143482
rect 324410 142488 324466 142497
rect 324410 142423 324466 142432
rect 324412 142112 324464 142118
rect 324412 142054 324464 142060
rect 324320 142044 324372 142050
rect 324320 141986 324372 141992
rect 324332 141681 324360 141986
rect 324318 141672 324374 141681
rect 324318 141607 324374 141616
rect 324424 140865 324452 142054
rect 324410 140856 324466 140865
rect 324410 140791 324466 140800
rect 324320 140752 324372 140758
rect 324320 140694 324372 140700
rect 324332 140185 324360 140694
rect 324318 140176 324374 140185
rect 324318 140111 324374 140120
rect 324412 139392 324464 139398
rect 324318 139360 324374 139369
rect 324412 139334 324464 139340
rect 324318 139295 324320 139304
rect 324372 139295 324374 139304
rect 324320 139266 324372 139272
rect 324424 138553 324452 139334
rect 324410 138544 324466 138553
rect 324410 138479 324466 138488
rect 324320 137964 324372 137970
rect 324320 137906 324372 137912
rect 324332 137873 324360 137906
rect 324412 137896 324464 137902
rect 324318 137864 324374 137873
rect 324412 137838 324464 137844
rect 324318 137799 324374 137808
rect 324424 137057 324452 137838
rect 324410 137048 324466 137057
rect 324410 136983 324466 136992
rect 324320 136604 324372 136610
rect 324320 136546 324372 136552
rect 324332 136377 324360 136546
rect 324318 136368 324374 136377
rect 324318 136303 324374 136312
rect 324964 136264 325016 136270
rect 324964 136206 325016 136212
rect 324320 135176 324372 135182
rect 324320 135118 324372 135124
rect 324332 134745 324360 135118
rect 324318 134736 324374 134745
rect 324318 134671 324374 134680
rect 324320 133884 324372 133890
rect 324320 133826 324372 133832
rect 324332 133249 324360 133826
rect 324318 133240 324374 133249
rect 324318 133175 324374 133184
rect 324412 132456 324464 132462
rect 324318 132424 324374 132433
rect 324412 132398 324464 132404
rect 324318 132359 324320 132368
rect 324372 132359 324374 132368
rect 324320 132330 324372 132336
rect 324424 131753 324452 132398
rect 324410 131744 324466 131753
rect 324410 131679 324466 131688
rect 324412 131096 324464 131102
rect 324412 131038 324464 131044
rect 324320 131028 324372 131034
rect 324320 130970 324372 130976
rect 324332 130937 324360 130970
rect 324318 130928 324374 130937
rect 324318 130863 324374 130872
rect 324424 130121 324452 131038
rect 324410 130112 324466 130121
rect 324410 130047 324466 130056
rect 324412 129736 324464 129742
rect 324412 129678 324464 129684
rect 324320 129668 324372 129674
rect 324320 129610 324372 129616
rect 324332 129441 324360 129610
rect 324318 129432 324374 129441
rect 324318 129367 324374 129376
rect 324424 128625 324452 129678
rect 324410 128616 324466 128625
rect 324410 128551 324466 128560
rect 324320 128308 324372 128314
rect 324320 128250 324372 128256
rect 324332 127809 324360 128250
rect 324318 127800 324374 127809
rect 324318 127735 324374 127744
rect 324320 126948 324372 126954
rect 324320 126890 324372 126896
rect 324332 126313 324360 126890
rect 324318 126304 324374 126313
rect 324318 126239 324374 126248
rect 324976 125497 325004 136206
rect 324962 125488 325018 125497
rect 324962 125423 325018 125432
rect 325606 124808 325662 124817
rect 325712 124794 325740 290527
rect 325804 134065 325832 299542
rect 329840 286340 329892 286346
rect 329840 286282 329892 286288
rect 328460 277500 328512 277506
rect 328460 277442 328512 277448
rect 327080 253972 327132 253978
rect 327080 253914 327132 253920
rect 325884 189780 325936 189786
rect 325884 189722 325936 189728
rect 325896 150929 325924 189722
rect 325974 175944 326030 175953
rect 325974 175879 326030 175888
rect 325988 171193 326016 175879
rect 325974 171184 326030 171193
rect 325974 171119 326030 171128
rect 325882 150920 325938 150929
rect 325882 150855 325938 150864
rect 327092 136270 327120 253914
rect 327172 250504 327224 250510
rect 327172 250446 327224 250452
rect 327184 150278 327212 250446
rect 327264 242208 327316 242214
rect 327264 242150 327316 242156
rect 327276 161906 327304 242150
rect 327356 185836 327408 185842
rect 327356 185778 327408 185784
rect 327264 161900 327316 161906
rect 327264 161842 327316 161848
rect 327368 153814 327396 185778
rect 327356 153808 327408 153814
rect 327356 153750 327408 153756
rect 327172 150272 327224 150278
rect 327172 150214 327224 150220
rect 327080 136264 327132 136270
rect 327080 136206 327132 136212
rect 325790 134056 325846 134065
rect 325790 133991 325846 134000
rect 328472 126954 328500 277442
rect 328552 231124 328604 231130
rect 328552 231066 328604 231072
rect 328564 128314 328592 231066
rect 328644 195288 328696 195294
rect 328644 195230 328696 195236
rect 328656 157350 328684 195230
rect 328734 178664 328790 178673
rect 328734 178599 328790 178608
rect 328644 157344 328696 157350
rect 328644 157286 328696 157292
rect 328748 146198 328776 178599
rect 328736 146192 328788 146198
rect 328736 146134 328788 146140
rect 329852 140758 329880 286282
rect 329932 271176 329984 271182
rect 329932 271118 329984 271124
rect 329944 144838 329972 271118
rect 331220 258120 331272 258126
rect 331220 258062 331272 258068
rect 330024 240168 330076 240174
rect 330024 240110 330076 240116
rect 329932 144832 329984 144838
rect 329932 144774 329984 144780
rect 329840 140752 329892 140758
rect 329840 140694 329892 140700
rect 330036 133890 330064 240110
rect 330116 218748 330168 218754
rect 330116 218690 330168 218696
rect 330024 133884 330076 133890
rect 330024 133826 330076 133832
rect 330128 129674 330156 218690
rect 331232 131034 331260 258062
rect 334072 221468 334124 221474
rect 334072 221410 334124 221416
rect 332876 206304 332928 206310
rect 332876 206246 332928 206252
rect 331312 186992 331364 186998
rect 331312 186934 331364 186940
rect 331324 139330 331352 186934
rect 331404 185632 331456 185638
rect 331404 185574 331456 185580
rect 331416 144906 331444 185574
rect 332692 181620 332744 181626
rect 332692 181562 332744 181568
rect 331496 178696 331548 178702
rect 331496 178638 331548 178644
rect 331508 162858 331536 178638
rect 332600 177540 332652 177546
rect 332600 177482 332652 177488
rect 332612 168298 332640 177482
rect 332600 168292 332652 168298
rect 332600 168234 332652 168240
rect 331496 162852 331548 162858
rect 331496 162794 331548 162800
rect 331404 144900 331456 144906
rect 331404 144842 331456 144848
rect 331312 139324 331364 139330
rect 331312 139266 331364 139272
rect 331220 131028 331272 131034
rect 331220 130970 331272 130976
rect 330116 129668 330168 129674
rect 330116 129610 330168 129616
rect 328552 128308 328604 128314
rect 328552 128250 328604 128256
rect 328460 126948 328512 126954
rect 328460 126890 328512 126896
rect 325662 124766 325740 124794
rect 325606 124743 325662 124752
rect 324320 124160 324372 124166
rect 324320 124102 324372 124108
rect 324332 123185 324360 124102
rect 324318 123176 324374 123185
rect 324318 123111 324374 123120
rect 324320 122800 324372 122806
rect 324320 122742 324372 122748
rect 324332 122505 324360 122742
rect 324318 122496 324374 122505
rect 324318 122431 324374 122440
rect 323122 121680 323178 121689
rect 323122 121615 323178 121624
rect 324412 121440 324464 121446
rect 324412 121382 324464 121388
rect 324320 121372 324372 121378
rect 324320 121314 324372 121320
rect 324332 120873 324360 121314
rect 324318 120864 324374 120873
rect 324318 120799 324374 120808
rect 324424 120193 324452 121382
rect 324410 120184 324466 120193
rect 324410 120119 324466 120128
rect 324320 120080 324372 120086
rect 324320 120022 324372 120028
rect 324332 119377 324360 120022
rect 324318 119368 324374 119377
rect 324318 119303 324374 119312
rect 324320 118652 324372 118658
rect 324320 118594 324372 118600
rect 324332 118561 324360 118594
rect 332704 118590 332732 181562
rect 332784 180192 332836 180198
rect 332784 180134 332836 180140
rect 332796 168366 332824 180134
rect 332784 168360 332836 168366
rect 332784 168302 332836 168308
rect 332888 139398 332916 206246
rect 333980 177404 334032 177410
rect 333980 177346 334032 177352
rect 332876 139392 332928 139398
rect 332876 139334 332928 139340
rect 324412 118584 324464 118590
rect 324318 118552 324374 118561
rect 324412 118526 324464 118532
rect 332692 118584 332744 118590
rect 332692 118526 332744 118532
rect 324318 118487 324374 118496
rect 324424 117881 324452 118526
rect 324410 117872 324466 117881
rect 324410 117807 324466 117816
rect 333992 117298 334020 177346
rect 334084 164150 334112 221410
rect 334636 194585 334664 302194
rect 345112 298240 345164 298246
rect 345112 298182 345164 298188
rect 335360 298172 335412 298178
rect 335360 298114 335412 298120
rect 334622 194576 334678 194585
rect 334622 194511 334678 194520
rect 334164 188556 334216 188562
rect 334164 188498 334216 188504
rect 334072 164144 334124 164150
rect 334072 164086 334124 164092
rect 334176 143478 334204 188498
rect 334256 185700 334308 185706
rect 334256 185642 334308 185648
rect 334268 150414 334296 185642
rect 334256 150408 334308 150414
rect 334256 150350 334308 150356
rect 335372 147626 335400 298114
rect 338120 296812 338172 296818
rect 338120 296754 338172 296760
rect 336740 295384 336792 295390
rect 336740 295326 336792 295332
rect 335452 207664 335504 207670
rect 335452 207606 335504 207612
rect 335360 147620 335412 147626
rect 335360 147562 335412 147568
rect 334164 143472 334216 143478
rect 334164 143414 334216 143420
rect 335464 137902 335492 207606
rect 335544 180124 335596 180130
rect 335544 180066 335596 180072
rect 335452 137896 335504 137902
rect 335452 137838 335504 137844
rect 324320 117292 324372 117298
rect 324320 117234 324372 117240
rect 333980 117292 334032 117298
rect 333980 117234 334032 117240
rect 324332 116385 324360 117234
rect 324318 116376 324374 116385
rect 324318 116311 324374 116320
rect 323490 115016 323546 115025
rect 323490 114951 323546 114960
rect 323504 114617 323532 114951
rect 323490 114608 323546 114617
rect 323490 114543 323546 114552
rect 324320 114504 324372 114510
rect 324320 114446 324372 114452
rect 324332 114073 324360 114446
rect 335556 114442 335584 180066
rect 335636 177472 335688 177478
rect 335636 177414 335688 177420
rect 335648 167006 335676 177414
rect 335636 167000 335688 167006
rect 335636 166942 335688 166948
rect 336752 122806 336780 295326
rect 336832 191208 336884 191214
rect 336832 191150 336884 191156
rect 336844 172514 336872 191150
rect 336924 182980 336976 182986
rect 336924 182922 336976 182928
rect 336832 172508 336884 172514
rect 336832 172450 336884 172456
rect 336936 158642 336964 182922
rect 337016 177336 337068 177342
rect 337016 177278 337068 177284
rect 336924 158636 336976 158642
rect 336924 158578 336976 158584
rect 336740 122800 336792 122806
rect 336740 122742 336792 122748
rect 324412 114436 324464 114442
rect 324412 114378 324464 114384
rect 335544 114436 335596 114442
rect 335544 114378 335596 114384
rect 324318 114064 324374 114073
rect 324318 113999 324374 114008
rect 324424 113257 324452 114378
rect 324410 113248 324466 113257
rect 324410 113183 324466 113192
rect 337028 113150 337056 177278
rect 338132 171086 338160 296754
rect 342904 296744 342956 296750
rect 342904 296686 342956 296692
rect 339498 295488 339554 295497
rect 339498 295423 339554 295432
rect 338396 199640 338448 199646
rect 338396 199582 338448 199588
rect 338212 184340 338264 184346
rect 338212 184282 338264 184288
rect 338120 171080 338172 171086
rect 338120 171022 338172 171028
rect 338224 120086 338252 184282
rect 338304 179376 338356 179382
rect 338302 179344 338304 179353
rect 338356 179344 338358 179353
rect 338302 179279 338358 179288
rect 338408 176050 338436 199582
rect 338488 182912 338540 182918
rect 338488 182854 338540 182860
rect 338396 176044 338448 176050
rect 338396 175986 338448 175992
rect 338500 175930 338528 182854
rect 338316 175902 338528 175930
rect 338316 121378 338344 175902
rect 338396 175840 338448 175846
rect 338396 175782 338448 175788
rect 338408 161362 338436 175782
rect 338396 161356 338448 161362
rect 338396 161298 338448 161304
rect 339512 135182 339540 295423
rect 342260 294024 342312 294030
rect 342260 293966 342312 293972
rect 340880 291304 340932 291310
rect 340878 291272 340880 291281
rect 340932 291272 340934 291281
rect 340878 291207 340934 291216
rect 339592 264988 339644 264994
rect 339592 264930 339644 264936
rect 339604 142050 339632 264930
rect 340880 262268 340932 262274
rect 340880 262210 340932 262216
rect 339776 203584 339828 203590
rect 339776 203526 339828 203532
rect 339684 181484 339736 181490
rect 339684 181426 339736 181432
rect 339592 142044 339644 142050
rect 339592 141986 339644 141992
rect 339500 135176 339552 135182
rect 339500 135118 339552 135124
rect 338304 121372 338356 121378
rect 338304 121314 338356 121320
rect 338212 120080 338264 120086
rect 338212 120022 338264 120028
rect 324320 113144 324372 113150
rect 324320 113086 324372 113092
rect 337016 113144 337068 113150
rect 337016 113086 337068 113092
rect 324332 112441 324360 113086
rect 324318 112432 324374 112441
rect 324318 112367 324374 112376
rect 323490 111208 323546 111217
rect 323490 111143 323546 111152
rect 323504 110537 323532 111143
rect 323490 110528 323546 110537
rect 323490 110463 323546 110472
rect 324320 108996 324372 109002
rect 324320 108938 324372 108944
rect 324332 108633 324360 108938
rect 324318 108624 324374 108633
rect 324318 108559 324374 108568
rect 324318 104816 324374 104825
rect 324318 104751 324374 104760
rect 323030 103184 323086 103193
rect 323030 103119 323086 103128
rect 324332 100314 324360 104751
rect 339696 103494 339724 181426
rect 339788 146266 339816 203526
rect 339776 146260 339828 146266
rect 339776 146202 339828 146208
rect 340892 124166 340920 262210
rect 340972 202156 341024 202162
rect 340972 202098 341024 202104
rect 340880 124160 340932 124166
rect 340880 124102 340932 124108
rect 340984 118658 341012 202098
rect 341062 182880 341118 182889
rect 341062 182815 341118 182824
rect 341076 136610 341104 182815
rect 341156 181552 341208 181558
rect 341156 181494 341208 181500
rect 341168 158710 341196 181494
rect 341156 158704 341208 158710
rect 341156 158646 341208 158652
rect 342272 142118 342300 293966
rect 342916 259418 342944 296686
rect 345020 282940 345072 282946
rect 345020 282882 345072 282888
rect 343732 266416 343784 266422
rect 343732 266358 343784 266364
rect 343640 260908 343692 260914
rect 343640 260850 343692 260856
rect 342904 259412 342956 259418
rect 342904 259354 342956 259360
rect 342352 224256 342404 224262
rect 342352 224198 342404 224204
rect 342260 142112 342312 142118
rect 342260 142054 342312 142060
rect 341064 136604 341116 136610
rect 341064 136546 341116 136552
rect 340972 118652 341024 118658
rect 340972 118594 341024 118600
rect 342364 114510 342392 224198
rect 342442 188320 342498 188329
rect 342442 188255 342498 188264
rect 342456 131102 342484 188255
rect 342536 181688 342588 181694
rect 342536 181630 342588 181636
rect 342548 153202 342576 181630
rect 342536 153196 342588 153202
rect 342536 153138 342588 153144
rect 343652 137970 343680 260850
rect 343744 149054 343772 266358
rect 343824 205012 343876 205018
rect 343824 204954 343876 204960
rect 343732 149048 343784 149054
rect 343732 148990 343784 148996
rect 343640 137964 343692 137970
rect 343640 137906 343692 137912
rect 342444 131096 342496 131102
rect 342444 131038 342496 131044
rect 343836 121446 343864 204954
rect 343916 191140 343968 191146
rect 343916 191082 343968 191088
rect 343928 165578 343956 191082
rect 343916 165572 343968 165578
rect 343916 165514 343968 165520
rect 345032 132394 345060 282882
rect 345124 161430 345152 298182
rect 346400 296880 346452 296886
rect 346400 296822 346452 296828
rect 345204 188352 345256 188358
rect 345204 188294 345256 188300
rect 345112 161424 345164 161430
rect 345112 161366 345164 161372
rect 345216 160070 345244 188294
rect 345296 182844 345348 182850
rect 345296 182786 345348 182792
rect 345308 164218 345336 182786
rect 345296 164212 345348 164218
rect 345296 164154 345348 164160
rect 345204 160064 345256 160070
rect 345204 160006 345256 160012
rect 346412 132462 346440 296822
rect 351920 287088 351972 287094
rect 351920 287030 351972 287036
rect 346492 277432 346544 277438
rect 346492 277374 346544 277380
rect 346504 155854 346532 277374
rect 347872 193928 347924 193934
rect 347872 193870 347924 193876
rect 347780 191276 347832 191282
rect 347780 191218 347832 191224
rect 346584 185904 346636 185910
rect 346584 185846 346636 185852
rect 346492 155848 346544 155854
rect 346492 155790 346544 155796
rect 346400 132456 346452 132462
rect 346400 132398 346452 132404
rect 345020 132388 345072 132394
rect 345020 132330 345072 132336
rect 346596 129742 346624 185846
rect 347792 151706 347820 191218
rect 347884 154562 347912 193870
rect 347964 193860 348016 193866
rect 347964 193802 348016 193808
rect 347976 155922 348004 193802
rect 347964 155916 348016 155922
rect 347964 155858 348016 155864
rect 347872 154556 347924 154562
rect 347872 154498 347924 154504
rect 347780 151700 347832 151706
rect 347780 151642 347832 151648
rect 351932 143546 351960 287030
rect 353300 248464 353352 248470
rect 353300 248406 353352 248412
rect 351920 143540 351972 143546
rect 351920 143482 351972 143488
rect 346584 129736 346636 129742
rect 346584 129678 346636 129684
rect 343824 121440 343876 121446
rect 343824 121382 343876 121388
rect 342352 114504 342404 114510
rect 342352 114446 342404 114452
rect 353312 109002 353340 248406
rect 359476 237386 359504 699654
rect 393964 275324 394016 275330
rect 393964 275266 394016 275272
rect 392582 269784 392638 269793
rect 392582 269719 392638 269728
rect 359464 237380 359516 237386
rect 359464 237322 359516 237328
rect 392596 126954 392624 269719
rect 393976 153202 394004 275266
rect 542372 231810 542400 702406
rect 580920 697241 580948 702442
rect 580906 697232 580962 697241
rect 580906 697167 580962 697176
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 582378 630864 582434 630873
rect 582378 630799 582434 630808
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 580262 325272 580318 325281
rect 580262 325207 580318 325216
rect 580276 312594 580304 325207
rect 580264 312588 580316 312594
rect 580264 312530 580316 312536
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580184 309806 580212 312015
rect 580172 309800 580224 309806
rect 580172 309742 580224 309748
rect 580262 289232 580318 289241
rect 580262 289167 580318 289176
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580184 271930 580212 272167
rect 580172 271924 580224 271930
rect 580172 271866 580224 271872
rect 579804 259412 579856 259418
rect 579804 259354 579856 259360
rect 579816 258913 579844 259354
rect 579802 258904 579858 258913
rect 579802 258839 579858 258848
rect 579894 245576 579950 245585
rect 579894 245511 579950 245520
rect 579908 244322 579936 245511
rect 579896 244316 579948 244322
rect 579896 244258 579948 244264
rect 542360 231804 542412 231810
rect 542360 231746 542412 231752
rect 574742 226944 574798 226953
rect 574742 226879 574798 226888
rect 574756 193186 574784 226879
rect 580172 206984 580224 206990
rect 580172 206926 580224 206932
rect 580184 205737 580212 206926
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 574744 193180 574796 193186
rect 574744 193122 574796 193128
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 393964 153196 394016 153202
rect 393964 153138 394016 153144
rect 579804 153196 579856 153202
rect 579804 153138 579856 153144
rect 579816 152697 579844 153138
rect 579802 152688 579858 152697
rect 579802 152623 579858 152632
rect 392584 126948 392636 126954
rect 392584 126890 392636 126896
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 353300 108996 353352 109002
rect 353300 108938 353352 108944
rect 324412 103488 324464 103494
rect 324412 103430 324464 103436
rect 339684 103488 339736 103494
rect 339684 103430 339736 103436
rect 324424 102513 324452 103430
rect 324410 102504 324466 102513
rect 324410 102439 324466 102448
rect 324332 100286 324452 100314
rect 324318 100192 324374 100201
rect 324318 100127 324374 100136
rect 324332 95198 324360 100127
rect 324320 95192 324372 95198
rect 324320 95134 324372 95140
rect 324424 95130 324452 100286
rect 324502 97064 324558 97073
rect 324502 96999 324558 97008
rect 324412 95124 324464 95130
rect 324412 95066 324464 95072
rect 321652 93832 321704 93838
rect 321652 93774 321704 93780
rect 324516 93770 324544 96999
rect 324504 93764 324556 93770
rect 324504 93706 324556 93712
rect 321560 93696 321612 93702
rect 321560 93638 321612 93644
rect 307300 91792 307352 91798
rect 307300 91734 307352 91740
rect 307208 90364 307260 90370
rect 307208 90306 307260 90312
rect 307116 89004 307168 89010
rect 307116 88946 307168 88952
rect 580276 73001 580304 289167
rect 580356 262880 580408 262886
rect 580356 262822 580408 262828
rect 580368 232393 580396 262822
rect 582392 257378 582420 630799
rect 582562 365120 582618 365129
rect 582562 365055 582618 365064
rect 582470 298208 582526 298217
rect 582470 298143 582526 298152
rect 582380 257372 582432 257378
rect 582380 257314 582432 257320
rect 582380 238060 582432 238066
rect 582380 238002 582432 238008
rect 580354 232384 580410 232393
rect 580354 232319 580410 232328
rect 580262 72992 580318 73001
rect 580262 72927 580318 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 307024 37936 307076 37942
rect 307024 37878 307076 37884
rect 305736 28348 305788 28354
rect 305736 28290 305788 28296
rect 305644 24200 305696 24206
rect 305644 24142 305696 24148
rect 304264 17332 304316 17338
rect 304264 17274 304316 17280
rect 298744 15972 298796 15978
rect 298744 15914 298796 15920
rect 297364 7676 297416 7682
rect 297364 7618 297416 7624
rect 582392 6633 582420 238002
rect 582484 19825 582512 298143
rect 582576 230450 582604 365055
rect 583024 299532 583076 299538
rect 583024 299474 583076 299480
rect 582654 298752 582710 298761
rect 582654 298687 582710 298696
rect 582668 234598 582696 298687
rect 582930 295352 582986 295361
rect 582930 295287 582986 295296
rect 582748 291236 582800 291242
rect 582748 291178 582800 291184
rect 582656 234592 582708 234598
rect 582656 234534 582708 234540
rect 582564 230444 582616 230450
rect 582564 230386 582616 230392
rect 582564 228404 582616 228410
rect 582564 228346 582616 228352
rect 582576 33153 582604 228346
rect 582760 112849 582788 291178
rect 582838 232520 582894 232529
rect 582838 232455 582894 232464
rect 582746 112840 582802 112849
rect 582746 112775 582802 112784
rect 582852 86193 582880 232455
rect 582944 179217 582972 295287
rect 583036 219065 583064 299474
rect 583116 235272 583168 235278
rect 583116 235214 583168 235220
rect 583022 219056 583078 219065
rect 583022 218991 583078 219000
rect 582930 179208 582986 179217
rect 582930 179143 582986 179152
rect 582838 86184 582894 86193
rect 582838 86119 582894 86128
rect 583128 46345 583156 235214
rect 583114 46336 583170 46345
rect 583114 46271 583170 46280
rect 582562 33144 582618 33153
rect 582562 33079 582618 33088
rect 582470 19816 582526 19825
rect 582470 19751 582526 19760
rect 582378 6624 582434 6633
rect 582378 6559 582434 6568
rect 295984 2100 296036 2106
rect 295984 2042 296036 2048
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3330 579944 3386 580000
rect 3238 566888 3294 566944
rect 3330 553832 3386 553888
rect 2962 527856 3018 527912
rect 3330 501744 3386 501800
rect 3054 475632 3110 475688
rect 3330 462576 3386 462632
rect 3330 449520 3386 449576
rect 2778 423564 2834 423600
rect 2778 423544 2780 423564
rect 2780 423544 2832 423564
rect 2832 423544 2834 423564
rect 3330 410488 3386 410544
rect 3330 397468 3332 397488
rect 3332 397468 3384 397488
rect 3384 397468 3386 397488
rect 3330 397432 3386 397468
rect 3330 371320 3386 371376
rect 3330 358400 3386 358456
rect 3330 345344 3386 345400
rect 3514 671200 3570 671256
rect 3514 658144 3570 658200
rect 3514 632068 3516 632088
rect 3516 632068 3568 632088
rect 3568 632068 3570 632088
rect 3514 632032 3570 632068
rect 3514 619112 3570 619168
rect 3514 606056 3570 606112
rect 3514 514800 3570 514856
rect 3330 319232 3386 319288
rect 3238 306176 3294 306232
rect 2778 293120 2834 293176
rect 3146 254088 3202 254144
rect 3054 241032 3110 241088
rect 3330 214920 3386 214976
rect 3054 201864 3110 201920
rect 3238 162832 3294 162888
rect 3146 110608 3202 110664
rect 2778 97552 2834 97608
rect 3606 267144 3662 267200
rect 3514 188808 3570 188864
rect 3514 149776 3570 149832
rect 3514 136720 3570 136776
rect 3514 84632 3570 84688
rect 3514 71576 3570 71632
rect 3422 58520 3478 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3146 32408 3202 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 6458 4800 6514 4856
rect 8298 61376 8354 61432
rect 15198 57160 15254 57216
rect 12438 54440 12494 54496
rect 11058 18536 11114 18592
rect 49606 210296 49662 210352
rect 50986 211792 51042 211848
rect 35898 62736 35954 62792
rect 49698 47504 49754 47560
rect 47582 32408 47638 32464
rect 59082 218592 59138 218648
rect 59266 179968 59322 180024
rect 75182 313928 75238 313984
rect 68650 300872 68706 300928
rect 67638 290536 67694 290592
rect 68834 296792 68890 296848
rect 68742 290128 68798 290184
rect 68650 289720 68706 289776
rect 68742 288768 68798 288824
rect 67730 287000 67786 287056
rect 67638 286728 67694 286784
rect 68282 285776 68338 285832
rect 67638 284688 67694 284744
rect 67638 283192 67694 283248
rect 67546 283056 67602 283112
rect 67362 280472 67418 280528
rect 64602 203496 64658 203552
rect 62026 190984 62082 191040
rect 67270 269456 67326 269512
rect 67638 280336 67694 280392
rect 67638 279112 67694 279168
rect 67730 278976 67786 279032
rect 67730 277752 67786 277808
rect 67638 277616 67694 277672
rect 67638 276392 67694 276448
rect 68006 276256 68062 276312
rect 67638 275032 67694 275088
rect 67730 274488 67786 274544
rect 68006 273536 68062 273592
rect 67730 272312 67786 272368
rect 67638 272176 67694 272232
rect 67638 270952 67694 271008
rect 67638 269592 67694 269648
rect 67638 268096 67694 268152
rect 67730 267416 67786 267472
rect 67638 267008 67694 267064
rect 67638 265376 67694 265432
rect 67730 264968 67786 265024
rect 67730 264152 67786 264208
rect 67638 263644 67640 263664
rect 67640 263644 67692 263664
rect 67692 263644 67694 263664
rect 67638 263608 67694 263644
rect 67638 263508 67640 263528
rect 67640 263508 67692 263528
rect 67692 263508 67694 263528
rect 67638 263472 67694 263508
rect 67638 262268 67694 262304
rect 67638 262248 67640 262268
rect 67640 262248 67692 262268
rect 67692 262248 67694 262268
rect 67730 261432 67786 261488
rect 67638 260924 67640 260944
rect 67640 260924 67692 260944
rect 67692 260924 67694 260944
rect 67638 260888 67694 260924
rect 67638 260788 67640 260808
rect 67640 260788 67692 260808
rect 67692 260788 67694 260808
rect 67638 260752 67694 260788
rect 67638 259528 67694 259584
rect 67730 258576 67786 258632
rect 67638 258188 67694 258224
rect 67638 258168 67640 258188
rect 67640 258168 67692 258188
rect 67692 258168 67694 258188
rect 68926 289448 68982 289504
rect 68834 288088 68890 288144
rect 68742 282104 68798 282160
rect 68374 275168 68430 275224
rect 67638 257216 67694 257272
rect 67638 255856 67694 255912
rect 67730 255332 67786 255368
rect 67730 255312 67732 255332
rect 67732 255312 67784 255332
rect 67784 255312 67786 255332
rect 67638 255212 67640 255232
rect 67640 255212 67692 255232
rect 67692 255212 67694 255232
rect 67638 255176 67694 255212
rect 67730 253136 67786 253192
rect 67638 252728 67694 252784
rect 67638 251776 67694 251832
rect 67730 250416 67786 250472
rect 67638 249892 67694 249928
rect 67638 249872 67640 249892
rect 67640 249872 67692 249892
rect 67692 249872 67694 249892
rect 67638 249756 67694 249792
rect 67638 249736 67640 249756
rect 67640 249736 67692 249756
rect 67692 249736 67694 249756
rect 75826 294208 75882 294264
rect 95790 294072 95846 294128
rect 104162 292576 104218 292632
rect 106094 298152 106150 298208
rect 105450 292712 105506 292768
rect 109958 295296 110014 295352
rect 108210 291896 108266 291952
rect 111798 295432 111854 295488
rect 113178 293936 113234 293992
rect 69754 291236 69810 291272
rect 69754 291216 69756 291236
rect 69756 291216 69808 291236
rect 69808 291216 69810 291236
rect 119802 290536 119858 290592
rect 69018 270816 69074 270872
rect 69202 268232 69258 268288
rect 69110 251232 69166 251288
rect 67454 240216 67510 240272
rect 67638 248512 67694 248568
rect 67638 247696 67694 247752
rect 67730 247152 67786 247208
rect 67638 246608 67694 246664
rect 67730 245928 67786 245984
rect 67638 245248 67694 245304
rect 67638 244568 67694 244624
rect 67730 243888 67786 243944
rect 67638 241848 67694 241904
rect 120078 268640 120134 268696
rect 120078 250960 120134 251016
rect 69662 244160 69718 244216
rect 119802 240896 119858 240952
rect 69110 196560 69166 196616
rect 71778 182824 71834 182880
rect 73250 225528 73306 225584
rect 79322 192480 79378 192536
rect 60646 178608 60702 178664
rect 84382 222808 84438 222864
rect 92478 188264 92534 188320
rect 99286 183640 99342 183696
rect 97538 177656 97594 177712
rect 99286 177656 99342 177712
rect 118974 239808 119030 239864
rect 114558 213152 114614 213208
rect 110694 179424 110750 179480
rect 106186 177656 106242 177712
rect 107566 177656 107622 177712
rect 114466 177656 114522 177712
rect 112994 177112 113050 177168
rect 110694 176976 110750 177032
rect 121550 291760 121606 291816
rect 121550 290400 121606 290456
rect 121550 289756 121552 289776
rect 121552 289756 121604 289776
rect 121604 289756 121606 289776
rect 121550 289720 121606 289756
rect 121550 288360 121606 288416
rect 121734 291080 121790 291136
rect 122010 289040 122066 289096
rect 121642 286320 121698 286376
rect 122102 287000 122158 287056
rect 122286 285640 122342 285696
rect 121550 284960 121606 285016
rect 121642 284280 121698 284336
rect 121458 282940 121514 282976
rect 121458 282920 121460 282940
rect 121460 282920 121512 282940
rect 121512 282920 121514 282940
rect 121458 281596 121460 281616
rect 121460 281596 121512 281616
rect 121512 281596 121514 281616
rect 121458 281560 121514 281596
rect 121458 280236 121460 280256
rect 121460 280236 121512 280256
rect 121512 280236 121514 280256
rect 121458 280200 121514 280236
rect 121458 278860 121514 278896
rect 121458 278840 121460 278860
rect 121460 278840 121512 278860
rect 121512 278840 121514 278860
rect 121458 277480 121514 277536
rect 121458 276800 121514 276856
rect 121458 274760 121514 274816
rect 121458 274080 121514 274136
rect 121458 273400 121514 273456
rect 121642 283600 121698 283656
rect 121642 282240 121698 282296
rect 121642 280880 121698 280936
rect 121642 279520 121698 279576
rect 121642 278160 121698 278216
rect 121642 276120 121698 276176
rect 121550 272720 121606 272776
rect 121550 271360 121606 271416
rect 121458 270000 121514 270056
rect 122102 275440 122158 275496
rect 121458 267960 121514 268016
rect 121550 267280 121606 267336
rect 121458 266600 121514 266656
rect 121550 265920 121606 265976
rect 121458 265240 121514 265296
rect 121642 264560 121698 264616
rect 122102 264152 122158 264208
rect 121550 263880 121606 263936
rect 121458 263200 121514 263256
rect 121458 262520 121514 262576
rect 121458 261840 121514 261896
rect 120262 261160 120318 261216
rect 121458 259800 121514 259856
rect 121458 259120 121514 259176
rect 121550 258440 121606 258496
rect 121550 257760 121606 257816
rect 121458 257080 121514 257136
rect 121458 256400 121514 256456
rect 121642 255720 121698 255776
rect 121550 255040 121606 255096
rect 121458 254360 121514 254416
rect 122102 253680 122158 253736
rect 121550 253000 121606 253056
rect 121458 252320 121514 252376
rect 121458 251640 121514 251696
rect 121550 250280 121606 250336
rect 121458 249600 121514 249656
rect 121458 248920 121514 248976
rect 121458 248240 121514 248296
rect 120170 247560 120226 247616
rect 121550 246880 121606 246936
rect 121550 245520 121606 245576
rect 121458 244840 121514 244896
rect 121642 244160 121698 244216
rect 121458 243480 121514 243536
rect 121458 242820 121514 242856
rect 121458 242800 121460 242820
rect 121460 242800 121512 242820
rect 121512 242800 121514 242820
rect 121550 242120 121606 242176
rect 121458 240760 121514 240816
rect 121550 240116 121552 240136
rect 121552 240116 121604 240136
rect 121604 240116 121606 240136
rect 121550 240080 121606 240116
rect 127714 292712 127770 292768
rect 142802 253136 142858 253192
rect 116950 177656 117006 177712
rect 118606 177656 118662 177712
rect 121366 177656 121422 177712
rect 123758 176976 123814 177032
rect 100666 176704 100722 176760
rect 103334 176704 103390 176760
rect 104622 176704 104678 176760
rect 108118 176724 108174 176760
rect 108118 176704 108120 176724
rect 108120 176704 108172 176724
rect 108172 176704 108174 176724
rect 109958 176704 110014 176760
rect 115846 176704 115902 176760
rect 129462 177656 129518 177712
rect 132406 177656 132462 177712
rect 133786 177656 133842 177712
rect 128082 176976 128138 177032
rect 124494 176740 124496 176760
rect 124496 176740 124548 176760
rect 124548 176740 124550 176760
rect 124494 176704 124550 176740
rect 126058 176704 126114 176760
rect 130750 176704 130806 176760
rect 134798 176704 134854 176760
rect 136086 176704 136142 176760
rect 148230 176704 148286 176760
rect 100758 175344 100814 175400
rect 121918 175344 121974 175400
rect 128174 175344 128230 175400
rect 158902 175344 158958 175400
rect 113178 174936 113234 174992
rect 119434 174936 119490 174992
rect 168010 171536 168066 171592
rect 177302 294208 177358 294264
rect 66166 129240 66222 129296
rect 65154 126248 65210 126304
rect 66074 125160 66130 125216
rect 65982 123528 66038 123584
rect 64786 122848 64842 122904
rect 65982 122848 66038 122904
rect 65982 122576 66038 122632
rect 65982 91024 66038 91080
rect 67546 128016 67602 128072
rect 67454 120808 67510 120864
rect 67362 102312 67418 102368
rect 66166 94832 66222 94888
rect 67638 100680 67694 100736
rect 67546 93744 67602 93800
rect 164882 95104 164938 95160
rect 111982 94696 112038 94752
rect 113730 94696 113786 94752
rect 129370 94696 129426 94752
rect 151634 94696 151690 94752
rect 118054 93608 118110 93664
rect 85670 93472 85726 93528
rect 107750 93472 107806 93528
rect 120630 93472 120686 93528
rect 110142 93200 110198 93256
rect 85118 92384 85174 92440
rect 91650 92384 91706 92440
rect 95054 92404 95110 92440
rect 95054 92384 95056 92404
rect 95056 92384 95108 92404
rect 95108 92384 95110 92404
rect 75826 91160 75882 91216
rect 90638 91704 90694 91760
rect 86866 91160 86922 91216
rect 88062 91160 88118 91216
rect 89626 91160 89682 91216
rect 106002 92384 106058 92440
rect 102690 91704 102746 91760
rect 100022 91568 100078 91624
rect 99286 91432 99342 91488
rect 97814 91296 97870 91352
rect 99102 91296 99158 91352
rect 93766 91160 93822 91216
rect 95146 91160 95202 91216
rect 96526 91160 96582 91216
rect 97906 91160 97962 91216
rect 97814 81368 97870 81424
rect 99194 91160 99250 91216
rect 99194 80008 99250 80064
rect 101862 91432 101918 91488
rect 100574 91160 100630 91216
rect 102046 91296 102102 91352
rect 101954 91160 102010 91216
rect 99286 78512 99342 78568
rect 104254 91160 104310 91216
rect 104806 91160 104862 91216
rect 107566 91296 107622 91352
rect 106186 91160 106242 91216
rect 107474 91160 107530 91216
rect 59358 30912 59414 30968
rect 54942 12960 54998 13016
rect 77390 29552 77446 29608
rect 108946 91160 109002 91216
rect 109590 91160 109646 91216
rect 115478 92420 115480 92440
rect 115480 92420 115532 92440
rect 115532 92420 115534 92440
rect 115478 92384 115534 92420
rect 116766 92384 116822 92440
rect 120538 92384 120594 92440
rect 161478 94424 161534 94480
rect 133142 93608 133198 93664
rect 110326 92248 110382 92304
rect 115386 91704 115442 91760
rect 111430 91296 111486 91352
rect 114374 91296 114430 91352
rect 111246 91160 111302 91216
rect 112350 91160 112406 91216
rect 114466 91160 114522 91216
rect 114374 88168 114430 88224
rect 115846 91160 115902 91216
rect 117134 91160 117190 91216
rect 118606 91160 118662 91216
rect 119986 91160 120042 91216
rect 125506 92384 125562 92440
rect 125966 92404 126022 92440
rect 125966 92384 125968 92404
rect 125968 92384 126020 92404
rect 126020 92384 126022 92404
rect 122838 91432 122894 91488
rect 122746 91296 122802 91352
rect 122654 91160 122710 91216
rect 123482 91160 123538 91216
rect 124126 91160 124182 91216
rect 125414 91160 125470 91216
rect 130750 92384 130806 92440
rect 151726 92384 151782 92440
rect 152094 92384 152150 92440
rect 136454 92112 136510 92168
rect 126702 91704 126758 91760
rect 126518 91160 126574 91216
rect 128266 91160 128322 91216
rect 132406 91160 132462 91216
rect 134614 91160 134670 91216
rect 126702 89664 126758 89720
rect 161478 91568 161534 91624
rect 151266 91432 151322 91488
rect 166906 115776 166962 115832
rect 166906 97960 166962 98016
rect 168010 111732 168012 111752
rect 168012 111732 168064 111752
rect 168064 111732 168066 111752
rect 168010 111696 168066 111732
rect 168102 110064 168158 110120
rect 168010 108704 168066 108760
rect 178682 177248 178738 177304
rect 177302 95104 177358 95160
rect 188342 294072 188398 294128
rect 186962 176840 187018 176896
rect 198002 185544 198058 185600
rect 213918 176160 213974 176216
rect 213918 175072 213974 175128
rect 214562 174664 214618 174720
rect 213918 173712 213974 173768
rect 214010 173304 214066 173360
rect 213274 172352 213330 172408
rect 213918 171944 213974 172000
rect 213918 170720 213974 170776
rect 214470 170856 214526 170912
rect 214010 169652 214066 169688
rect 214010 169632 214012 169652
rect 214012 169632 214064 169652
rect 214064 169632 214066 169652
rect 213918 169360 213974 169416
rect 213918 168000 213974 168056
rect 214010 167864 214066 167920
rect 214470 166640 214526 166696
rect 213918 166096 213974 166152
rect 213918 165280 213974 165336
rect 214010 164736 214066 164792
rect 213918 164092 213920 164112
rect 213920 164092 213972 164112
rect 213972 164092 213974 164112
rect 213918 164056 213974 164092
rect 214010 163376 214066 163432
rect 213918 161472 213974 161528
rect 213918 161200 213974 161256
rect 214010 160792 214066 160848
rect 213918 160012 213920 160032
rect 213920 160012 213972 160032
rect 213972 160012 213974 160032
rect 213918 159976 213974 160012
rect 213918 158652 213920 158672
rect 213920 158652 213972 158672
rect 213972 158652 213974 158672
rect 213918 158616 213974 158652
rect 214010 158072 214066 158128
rect 213918 157276 213974 157312
rect 213918 157256 213920 157276
rect 213920 157256 213972 157276
rect 213972 157256 213974 157276
rect 214010 156848 214066 156904
rect 213918 155488 213974 155544
rect 214010 153856 214066 153912
rect 213918 153448 213974 153504
rect 213182 152632 213238 152688
rect 199382 94424 199438 94480
rect 207754 94832 207810 94888
rect 214378 152088 214434 152144
rect 213918 151952 213974 152008
rect 214010 150864 214066 150920
rect 213918 150048 213974 150104
rect 214746 166912 214802 166968
rect 214654 159432 214710 159488
rect 214654 150728 214710 150784
rect 214562 149504 214618 149560
rect 213918 148688 213974 148744
rect 213918 148008 213974 148064
rect 214010 146648 214066 146704
rect 213918 146376 213974 146432
rect 214010 145288 214066 145344
rect 213918 144916 213920 144936
rect 213920 144916 213972 144936
rect 213972 144916 213974 144936
rect 213918 144880 213974 144916
rect 214010 143928 214066 143984
rect 213918 143520 213974 143576
rect 213918 142180 213974 142216
rect 213918 142160 213920 142180
rect 213920 142160 213972 142180
rect 213972 142160 213974 142180
rect 214010 141344 214066 141400
rect 213918 140936 213974 140992
rect 214010 139984 214066 140040
rect 213918 139576 213974 139632
rect 214470 138760 214526 138816
rect 213918 138080 213974 138136
rect 213918 136720 213974 136776
rect 214010 135632 214066 135688
rect 213918 135360 213974 135416
rect 214010 134272 214066 134328
rect 213918 134020 213974 134056
rect 213918 134000 213920 134020
rect 213920 134000 213972 134020
rect 213972 134000 213974 134020
rect 214010 132776 214066 132832
rect 213918 132524 213974 132560
rect 213918 132504 213920 132524
rect 213920 132504 213972 132524
rect 213972 132504 213974 132524
rect 214654 137400 214710 137456
rect 214010 131416 214066 131472
rect 213918 131180 213920 131200
rect 213920 131180 213972 131200
rect 213972 131180 213974 131200
rect 213918 131144 213974 131180
rect 214010 130056 214066 130112
rect 213918 129804 213974 129840
rect 213918 129784 213920 129804
rect 213920 129784 213972 129804
rect 213972 129784 213974 129804
rect 213918 128832 213974 128888
rect 213458 127472 213514 127528
rect 213458 127064 213514 127120
rect 214010 126112 214066 126168
rect 213918 125704 213974 125760
rect 214010 124752 214066 124808
rect 213918 124344 213974 124400
rect 213918 123528 213974 123584
rect 213918 122868 213974 122904
rect 213918 122848 213920 122868
rect 213920 122848 213972 122868
rect 213972 122848 213974 122868
rect 214010 122168 214066 122224
rect 213918 121760 213974 121816
rect 213918 120808 213974 120864
rect 213274 120128 213330 120184
rect 214010 119584 214066 119640
rect 213918 118904 213974 118960
rect 214102 119040 214158 119096
rect 213366 117544 213422 117600
rect 213918 117308 213920 117328
rect 213920 117308 213972 117328
rect 213972 117308 213974 117328
rect 213918 117272 213974 117308
rect 214010 116184 214066 116240
rect 213918 115912 213974 115968
rect 214010 114960 214066 115016
rect 213918 114588 213920 114608
rect 213920 114588 213972 114608
rect 213972 114588 213974 114608
rect 213918 114552 213974 114588
rect 213918 113600 213974 113656
rect 214010 113228 214012 113248
rect 214012 113228 214064 113248
rect 214064 113228 214066 113248
rect 214010 113192 214066 113228
rect 214010 112240 214066 112296
rect 213918 111852 213974 111888
rect 213918 111832 213920 111852
rect 213920 111832 213972 111852
rect 213972 111832 213974 111852
rect 214010 110880 214066 110936
rect 213918 110492 213974 110528
rect 213918 110472 213920 110492
rect 213920 110472 213972 110492
rect 213972 110472 213974 110492
rect 214010 109656 214066 109712
rect 213918 109248 213974 109304
rect 213918 107888 213974 107944
rect 213918 106936 213974 106992
rect 214010 105712 214066 105768
rect 213918 105304 213974 105360
rect 213918 103944 213974 104000
rect 213918 103672 213974 103728
rect 214838 108296 214894 108352
rect 214654 106256 214710 106312
rect 214010 99728 214066 99784
rect 213918 99476 213974 99512
rect 213918 99456 213920 99476
rect 213920 99456 213972 99476
rect 213972 99456 213974 99476
rect 214010 98368 214066 98424
rect 213918 97996 213920 98016
rect 213920 97996 213972 98016
rect 213972 97996 213974 98016
rect 213918 97960 213974 97996
rect 214562 101088 214618 101144
rect 214470 97144 214526 97200
rect 213918 97008 213974 97064
rect 213918 95784 213974 95840
rect 214930 96600 214986 96656
rect 232502 177520 232558 177576
rect 226982 177384 227038 177440
rect 224222 176024 224278 176080
rect 245014 178744 245070 178800
rect 220082 175888 220138 175944
rect 246946 175752 247002 175808
rect 249246 175208 249302 175264
rect 249154 174664 249210 174720
rect 249154 172744 249210 172800
rect 217322 155352 217378 155408
rect 217322 154672 217378 154728
rect 249890 165688 249946 165744
rect 251178 158752 251234 158808
rect 249890 158208 249946 158264
rect 250442 155216 250498 155272
rect 249798 150728 249854 150784
rect 252466 173712 252522 173768
rect 252374 172352 252430 172408
rect 252466 171400 252522 171456
rect 252466 170176 252522 170232
rect 252466 170040 252522 170096
rect 252466 169496 252522 169552
rect 252374 169088 252430 169144
rect 252282 168544 252338 168600
rect 252282 167592 252338 167648
rect 252466 168136 252522 168192
rect 252374 167184 252430 167240
rect 252466 166640 252522 166696
rect 252374 166232 252430 166288
rect 252466 165280 252522 165336
rect 252374 164736 252430 164792
rect 252466 163920 252522 163976
rect 251454 162968 251510 163024
rect 252466 162424 252522 162480
rect 252374 162016 252430 162072
rect 252282 161472 252338 161528
rect 252466 160520 252522 160576
rect 251362 160112 251418 160168
rect 252466 159568 252522 159624
rect 252006 159160 252062 159216
rect 252466 157292 252468 157312
rect 252468 157292 252520 157312
rect 252520 157292 252522 157312
rect 252466 157256 252522 157292
rect 252466 156848 252522 156904
rect 252374 156304 252430 156360
rect 252466 155896 252522 155952
rect 251454 155352 251510 155408
rect 252374 154944 252430 155000
rect 252466 154436 252468 154456
rect 252468 154436 252520 154456
rect 252520 154436 252522 154456
rect 252466 154400 252522 154436
rect 252374 153992 252430 154048
rect 252466 153076 252468 153096
rect 252468 153076 252520 153096
rect 252520 153076 252522 153096
rect 252466 153040 252522 153076
rect 252650 171808 252706 171864
rect 252742 164328 252798 164384
rect 252558 152632 252614 152688
rect 252282 152088 252338 152144
rect 251270 146920 251326 146976
rect 250442 143656 250498 143712
rect 252466 151716 252468 151736
rect 252468 151716 252520 151736
rect 252520 151716 252522 151736
rect 252466 151680 252522 151716
rect 252006 151136 252062 151192
rect 252282 150220 252284 150240
rect 252284 150220 252336 150240
rect 252336 150220 252338 150240
rect 252282 150184 252338 150220
rect 252466 149776 252522 149832
rect 252374 149232 252430 149288
rect 252834 148824 252890 148880
rect 252466 148280 252522 148336
rect 252374 147872 252430 147928
rect 252466 146512 252522 146568
rect 252190 146240 252246 146296
rect 251362 140800 251418 140856
rect 216218 102448 216274 102504
rect 216126 100816 216182 100872
rect 249154 96600 249210 96656
rect 252466 145968 252522 146024
rect 252374 145560 252430 145616
rect 252282 145016 252338 145072
rect 252466 144064 252522 144120
rect 252190 142704 252246 142760
rect 252466 143112 252522 143168
rect 252374 142160 252430 142216
rect 252466 141344 252522 141400
rect 252466 139848 252522 139904
rect 252374 139440 252430 139496
rect 252006 136176 252062 136232
rect 252282 138488 252338 138544
rect 252374 137944 252430 138000
rect 252466 137536 252522 137592
rect 252282 136992 252338 137048
rect 252466 136584 252522 136640
rect 252282 135632 252338 135688
rect 252374 135224 252430 135280
rect 252466 134680 252522 134736
rect 252374 134272 252430 134328
rect 252466 133764 252468 133784
rect 252468 133764 252520 133784
rect 252520 133764 252522 133784
rect 252466 133728 252522 133764
rect 252374 133320 252430 133376
rect 252190 132776 252246 132832
rect 252374 132368 252430 132424
rect 252466 131824 252522 131880
rect 252282 131416 252338 131472
rect 252466 130464 252522 130520
rect 252282 130056 252338 130112
rect 251914 126248 251970 126304
rect 251638 117272 251694 117328
rect 252374 129512 252430 129568
rect 252466 129104 252522 129160
rect 252282 128560 252338 128616
rect 252466 128188 252468 128208
rect 252468 128188 252520 128208
rect 252520 128188 252522 128208
rect 252466 128152 252522 128188
rect 252374 127608 252430 127664
rect 252466 127200 252522 127256
rect 252466 126656 252522 126712
rect 252374 125704 252430 125760
rect 252374 125296 252430 125352
rect 252190 124344 252246 124400
rect 252466 124752 252522 124808
rect 252282 123936 252338 123992
rect 252466 123392 252522 123448
rect 252374 122984 252430 123040
rect 252466 122440 252522 122496
rect 253202 122032 253258 122088
rect 252374 121488 252430 121544
rect 252466 121080 252522 121136
rect 252374 120536 252430 120592
rect 252282 120128 252338 120184
rect 252466 119584 252522 119640
rect 252466 119176 252522 119232
rect 252374 118768 252430 118824
rect 252006 116864 252062 116920
rect 251914 110744 251970 110800
rect 251638 109792 251694 109848
rect 251178 103128 251234 103184
rect 252466 118224 252522 118280
rect 252374 117816 252430 117872
rect 252466 116320 252522 116376
rect 252466 115912 252522 115968
rect 252282 115368 252338 115424
rect 252374 114960 252430 115016
rect 252466 114452 252468 114472
rect 252468 114452 252520 114472
rect 252520 114452 252522 114472
rect 252466 114416 252522 114452
rect 252374 114008 252430 114064
rect 252282 113464 252338 113520
rect 252466 112104 252522 112160
rect 252374 111716 252430 111752
rect 252374 111696 252376 111716
rect 252376 111696 252428 111716
rect 252428 111696 252430 111716
rect 252466 111152 252522 111208
rect 252098 108840 252154 108896
rect 252466 110200 252522 110256
rect 252374 109248 252430 109304
rect 252466 108296 252522 108352
rect 252374 107888 252430 107944
rect 252282 106936 252338 106992
rect 252466 107516 252468 107536
rect 252468 107516 252520 107536
rect 252520 107516 252522 107536
rect 252466 107480 252522 107516
rect 252374 106528 252430 106584
rect 252466 105984 252522 106040
rect 252282 105576 252338 105632
rect 252190 105032 252246 105088
rect 252282 104080 252338 104136
rect 252006 103672 252062 103728
rect 252466 104624 252522 104680
rect 251362 101768 251418 101824
rect 252374 102720 252430 102776
rect 252466 102176 252522 102232
rect 252190 100816 252246 100872
rect 252466 101360 252522 101416
rect 252282 100408 252338 100464
rect 252466 99864 252522 99920
rect 252374 99456 252430 99512
rect 251270 98504 251326 98560
rect 252466 98912 252522 98968
rect 252374 97960 252430 98016
rect 252466 97552 252522 97608
rect 251270 97008 251326 97064
rect 252466 97008 252522 97064
rect 251178 96192 251234 96248
rect 252466 96600 252522 96656
rect 258998 142296 259054 142352
rect 300122 700304 300178 700360
rect 265622 145560 265678 145616
rect 332506 702480 332562 702536
rect 302882 178880 302938 178936
rect 298742 178744 298798 178800
rect 286322 177248 286378 177304
rect 307114 175208 307170 175264
rect 306562 174800 306618 174856
rect 306562 172216 306618 172272
rect 306562 170584 306618 170640
rect 307022 165008 307078 165064
rect 303526 148280 303582 148336
rect 306562 159024 306618 159080
rect 306930 158208 306986 158264
rect 305734 157392 305790 157448
rect 305642 145016 305698 145072
rect 306562 154808 306618 154864
rect 306562 154400 306618 154456
rect 306654 153176 306710 153232
rect 306930 151000 306986 151056
rect 306562 148824 306618 148880
rect 305918 147872 305974 147928
rect 305826 118768 305882 118824
rect 305642 110608 305698 110664
rect 305734 106664 305790 106720
rect 306930 146784 306986 146840
rect 306562 143384 306618 143440
rect 306562 142024 306618 142080
rect 306746 140800 306802 140856
rect 306562 139032 306618 139088
rect 306562 136176 306618 136232
rect 306930 139984 306986 140040
rect 307574 174392 307630 174448
rect 307666 174004 307722 174040
rect 307666 173984 307668 174004
rect 307668 173984 307720 174004
rect 307720 173984 307722 174004
rect 307574 173576 307630 173632
rect 307482 172660 307484 172680
rect 307484 172660 307536 172680
rect 307536 172660 307538 172680
rect 307482 172624 307538 172660
rect 307666 173168 307722 173224
rect 307574 171808 307630 171864
rect 307666 171400 307722 171456
rect 307574 170992 307630 171048
rect 307666 170176 307722 170232
rect 307390 169768 307446 169824
rect 307298 166368 307354 166424
rect 307298 165416 307354 165472
rect 307666 169224 307722 169280
rect 307574 168816 307630 168872
rect 307482 168444 307484 168464
rect 307484 168444 307536 168464
rect 307536 168444 307538 168464
rect 307482 168408 307538 168444
rect 307482 168000 307538 168056
rect 307574 167592 307630 167648
rect 307666 167204 307722 167240
rect 307666 167184 307668 167204
rect 307668 167184 307720 167204
rect 307720 167184 307722 167204
rect 307574 166776 307630 166832
rect 307666 165824 307722 165880
rect 307666 164600 307722 164656
rect 307574 164192 307630 164248
rect 307574 163784 307630 163840
rect 307482 163376 307538 163432
rect 307666 162968 307722 163024
rect 307574 162424 307630 162480
rect 307482 162016 307538 162072
rect 307666 161608 307722 161664
rect 307206 160792 307262 160848
rect 307574 161200 307630 161256
rect 307666 160384 307722 160440
rect 307298 159976 307354 160032
rect 307666 159568 307722 159624
rect 307574 158616 307630 158672
rect 307666 157800 307722 157856
rect 307482 156984 307538 157040
rect 307574 156576 307630 156632
rect 307666 156168 307722 156224
rect 307298 155624 307354 155680
rect 307666 155216 307722 155272
rect 307666 153584 307722 153640
rect 307482 152632 307538 152688
rect 307574 152224 307630 152280
rect 307666 151852 307668 151872
rect 307668 151852 307720 151872
rect 307720 151852 307722 151872
rect 307666 151816 307722 151852
rect 307298 151408 307354 151464
rect 307666 150612 307722 150648
rect 307666 150592 307668 150612
rect 307668 150592 307720 150612
rect 307720 150592 307722 150612
rect 307666 150184 307722 150240
rect 307390 149776 307446 149832
rect 307298 147192 307354 147248
rect 307114 145832 307170 145888
rect 307574 149232 307630 149288
rect 307482 147600 307538 147656
rect 307666 148416 307722 148472
rect 307390 144880 307446 144936
rect 307482 144608 307538 144664
rect 307574 144200 307630 144256
rect 307666 143792 307722 143848
rect 307206 140392 307262 140448
rect 307114 137808 307170 137864
rect 306746 128832 306802 128888
rect 306930 125024 306986 125080
rect 306562 118632 306618 118688
rect 306746 116592 306802 116648
rect 306010 107616 306066 107672
rect 306930 102992 306986 103048
rect 307022 98640 307078 98696
rect 306930 96600 306986 96656
rect 307298 139576 307354 139632
rect 307298 135632 307354 135688
rect 307206 132640 307262 132696
rect 307574 142976 307630 143032
rect 307666 142432 307722 142488
rect 307574 141616 307630 141672
rect 307666 141208 307722 141264
rect 307574 138624 307630 138680
rect 307666 138216 307722 138272
rect 307574 137400 307630 137456
rect 307666 136992 307722 137048
rect 307482 136584 307538 136640
rect 307666 135260 307668 135280
rect 307668 135260 307720 135280
rect 307720 135260 307722 135280
rect 307666 135224 307722 135260
rect 307390 132232 307446 132288
rect 307574 134816 307630 134872
rect 307666 134408 307722 134464
rect 307574 133592 307630 133648
rect 307666 133184 307722 133240
rect 307574 131824 307630 131880
rect 307666 131416 307722 131472
rect 307666 131008 307722 131064
rect 307298 124616 307354 124672
rect 307574 129920 307630 129976
rect 307482 129820 307484 129840
rect 307484 129820 307536 129840
rect 307536 129820 307538 129840
rect 307482 129784 307538 129820
rect 307574 129240 307630 129296
rect 307666 128444 307722 128480
rect 307666 128424 307668 128444
rect 307668 128424 307720 128444
rect 307720 128424 307722 128444
rect 307482 128016 307538 128072
rect 307574 127608 307630 127664
rect 307666 127200 307722 127256
rect 307482 126792 307538 126848
rect 307574 126384 307630 126440
rect 307666 125840 307722 125896
rect 307574 125432 307630 125488
rect 307666 124228 307722 124264
rect 307666 124208 307668 124228
rect 307668 124208 307720 124228
rect 307720 124208 307722 124228
rect 307482 123800 307538 123856
rect 307666 123392 307722 123448
rect 307574 122984 307630 123040
rect 307482 122440 307538 122496
rect 307574 122032 307630 122088
rect 307666 121624 307722 121680
rect 307482 121216 307538 121272
rect 307574 120808 307630 120864
rect 307666 120400 307722 120456
rect 307482 119992 307538 120048
rect 307574 119584 307630 119640
rect 307666 119040 307722 119096
rect 307574 118768 307630 118824
rect 307574 117816 307630 117872
rect 307666 117444 307668 117464
rect 307668 117444 307720 117464
rect 307720 117444 307722 117464
rect 307666 117408 307722 117444
rect 307574 117000 307630 117056
rect 307666 116184 307722 116240
rect 307482 115640 307538 115696
rect 307574 115232 307630 115288
rect 307666 114824 307722 114880
rect 307666 113600 307722 113656
rect 307574 113212 307630 113248
rect 307574 113192 307576 113212
rect 307576 113192 307628 113212
rect 307628 113192 307630 113212
rect 307666 111968 307722 112024
rect 307482 111868 307484 111888
rect 307484 111868 307536 111888
rect 307536 111868 307538 111888
rect 307482 111832 307538 111868
rect 307574 111424 307630 111480
rect 307666 111016 307722 111072
rect 307482 110200 307538 110256
rect 307574 109792 307630 109848
rect 307666 109248 307722 109304
rect 307482 108840 307538 108896
rect 307666 108432 307722 108488
rect 307574 108024 307630 108080
rect 307482 107616 307538 107672
rect 307666 107616 307722 107672
rect 307666 107208 307722 107264
rect 307482 106428 307484 106448
rect 307484 106428 307536 106448
rect 307536 106428 307538 106448
rect 307482 106392 307538 106428
rect 307482 105848 307538 105904
rect 307666 105440 307722 105496
rect 307574 105032 307630 105088
rect 307574 104624 307630 104680
rect 307666 103808 307722 103864
rect 307574 103400 307630 103456
rect 307666 102448 307722 102504
rect 307482 101632 307538 101688
rect 307574 101224 307630 101280
rect 307666 100816 307722 100872
rect 307574 100408 307630 100464
rect 307666 100000 307722 100056
rect 307574 99048 307630 99104
rect 307666 98232 307722 98288
rect 307666 97416 307722 97472
rect 307666 96192 307722 96248
rect 322938 292576 322994 292632
rect 309138 114416 309194 114472
rect 309138 113056 309194 113112
rect 316038 176704 316094 176760
rect 316314 176160 316370 176216
rect 321466 176024 321522 176080
rect 321466 175208 321522 175264
rect 321282 169632 321338 169688
rect 325698 290536 325754 290592
rect 322938 156984 322994 157040
rect 321742 148280 321798 148336
rect 321650 127472 321706 127528
rect 321558 124208 321614 124264
rect 321558 105032 321614 105088
rect 321282 98776 321338 98832
rect 321374 97280 321430 97336
rect 321282 95104 321338 95160
rect 321466 96620 321522 96656
rect 321466 96600 321468 96620
rect 321468 96600 321520 96620
rect 321520 96600 321522 96620
rect 321650 103672 321706 103728
rect 324318 172352 324374 172408
rect 324318 170856 324374 170912
rect 324502 173984 324558 174040
rect 324594 173168 324650 173224
rect 324410 168544 324466 168600
rect 324318 167728 324374 167784
rect 324410 167048 324466 167104
rect 324318 166232 324374 166288
rect 323214 165416 323270 165472
rect 324318 164736 324374 164792
rect 324318 163920 324374 163976
rect 324410 163104 324466 163160
rect 324318 162424 324374 162480
rect 324318 161608 324374 161664
rect 324318 160792 324374 160848
rect 324410 160112 324466 160168
rect 324318 159296 324374 159352
rect 324318 158480 324374 158536
rect 324410 157800 324466 157856
rect 324318 156304 324374 156360
rect 324318 155488 324374 155544
rect 324410 154672 324466 154728
rect 324318 153992 324374 154048
rect 324318 153176 324374 153232
rect 324410 152360 324466 152416
rect 324318 151700 324374 151736
rect 324318 151680 324320 151700
rect 324320 151680 324372 151700
rect 324372 151680 324374 151700
rect 324318 150048 324374 150104
rect 324410 149368 324466 149424
rect 324318 148552 324374 148608
rect 324318 147056 324374 147112
rect 324318 146260 324374 146296
rect 324318 146240 324320 146260
rect 324320 146240 324372 146260
rect 324372 146240 324374 146260
rect 324410 145424 324466 145480
rect 324318 144744 324374 144800
rect 324410 143928 324466 143984
rect 324318 143112 324374 143168
rect 324410 142432 324466 142488
rect 324318 141616 324374 141672
rect 324410 140800 324466 140856
rect 324318 140120 324374 140176
rect 324318 139324 324374 139360
rect 324318 139304 324320 139324
rect 324320 139304 324372 139324
rect 324372 139304 324374 139324
rect 324410 138488 324466 138544
rect 324318 137808 324374 137864
rect 324410 136992 324466 137048
rect 324318 136312 324374 136368
rect 324318 134680 324374 134736
rect 324318 133184 324374 133240
rect 324318 132388 324374 132424
rect 324318 132368 324320 132388
rect 324320 132368 324372 132388
rect 324372 132368 324374 132388
rect 324410 131688 324466 131744
rect 324318 130872 324374 130928
rect 324410 130056 324466 130112
rect 324318 129376 324374 129432
rect 324410 128560 324466 128616
rect 324318 127744 324374 127800
rect 324318 126248 324374 126304
rect 324962 125432 325018 125488
rect 325606 124752 325662 124808
rect 325974 175888 326030 175944
rect 325974 171128 326030 171184
rect 325882 150864 325938 150920
rect 325790 134000 325846 134056
rect 328734 178608 328790 178664
rect 324318 123120 324374 123176
rect 324318 122440 324374 122496
rect 323122 121624 323178 121680
rect 324318 120808 324374 120864
rect 324410 120128 324466 120184
rect 324318 119312 324374 119368
rect 324318 118496 324374 118552
rect 324410 117816 324466 117872
rect 334622 194520 334678 194576
rect 324318 116320 324374 116376
rect 323490 114960 323546 115016
rect 323490 114552 323546 114608
rect 324318 114008 324374 114064
rect 324410 113192 324466 113248
rect 339498 295432 339554 295488
rect 338302 179324 338304 179344
rect 338304 179324 338356 179344
rect 338356 179324 338358 179344
rect 338302 179288 338358 179324
rect 340878 291252 340880 291272
rect 340880 291252 340932 291272
rect 340932 291252 340934 291272
rect 340878 291216 340934 291252
rect 324318 112376 324374 112432
rect 323490 111152 323546 111208
rect 323490 110472 323546 110528
rect 324318 108568 324374 108624
rect 324318 104760 324374 104816
rect 323030 103128 323086 103184
rect 341062 182824 341118 182880
rect 342442 188264 342498 188320
rect 392582 269728 392638 269784
rect 580906 697176 580962 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 582378 630808 582434 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 431568 580226 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 580262 325216 580318 325272
rect 580170 312024 580226 312080
rect 580262 289176 580318 289232
rect 580170 272176 580226 272232
rect 579802 258848 579858 258904
rect 579894 245520 579950 245576
rect 574742 226888 574798 226944
rect 580170 205672 580226 205728
rect 580170 192480 580226 192536
rect 579802 152632 579858 152688
rect 580170 125976 580226 126032
rect 324410 102448 324466 102504
rect 324318 100136 324374 100192
rect 324502 97008 324558 97064
rect 582562 365064 582618 365120
rect 582470 298152 582526 298208
rect 580354 232328 580410 232384
rect 580262 72936 580318 72992
rect 580170 59608 580226 59664
rect 582654 298696 582710 298752
rect 582930 295296 582986 295352
rect 582838 232464 582894 232520
rect 582746 112784 582802 112840
rect 583022 219000 583078 219056
rect 582930 179152 582986 179208
rect 582838 86128 582894 86184
rect 583114 46280 583170 46336
rect 582562 33088 582618 33144
rect 582470 19760 582526 19816
rect 582378 6568 582434 6624
<< metal3 >>
rect 70894 702476 70900 702540
rect 70964 702538 70970 702540
rect 332501 702538 332567 702541
rect 70964 702536 332567 702538
rect 70964 702480 332506 702536
rect 332562 702480 332567 702536
rect 70964 702478 332567 702480
rect 70964 702476 70970 702478
rect 332501 702475 332567 702478
rect 59118 700300 59124 700364
rect 59188 700362 59194 700364
rect 300117 700362 300183 700365
rect 59188 700360 300183 700362
rect 59188 700304 300122 700360
rect 300178 700304 300183 700360
rect 59188 700302 300183 700304
rect 59188 700300 59194 700302
rect 300117 700299 300183 700302
rect -960 697220 480 697460
rect 580901 697234 580967 697237
rect 583520 697234 584960 697324
rect 580901 697232 584960 697234
rect 580901 697176 580906 697232
rect 580962 697176 584960 697232
rect 580901 697174 584960 697176
rect 580901 697171 580967 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 582373 630866 582439 630869
rect 583520 630866 584960 630956
rect 582373 630864 584960 630866
rect 582373 630808 582378 630864
rect 582434 630808 584960 630864
rect 582373 630806 584960 630808
rect 582373 630803 582439 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3233 566946 3299 566949
rect -960 566944 3299 566946
rect -960 566888 3238 566944
rect 3294 566888 3299 566944
rect -960 566886 3299 566888
rect -960 566796 480 566886
rect 3233 566883 3299 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3325 501802 3391 501805
rect -960 501800 3391 501802
rect -960 501744 3330 501800
rect 3386 501744 3391 501800
rect -960 501742 3391 501744
rect -960 501652 480 501742
rect 3325 501739 3391 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3049 475690 3115 475693
rect -960 475688 3115 475690
rect -960 475632 3054 475688
rect 3110 475632 3115 475688
rect -960 475630 3115 475632
rect -960 475540 480 475630
rect 3049 475627 3115 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3325 462634 3391 462637
rect -960 462632 3391 462634
rect -960 462576 3330 462632
rect 3386 462576 3391 462632
rect -960 462574 3391 462576
rect -960 462484 480 462574
rect 3325 462571 3391 462574
rect 583520 458146 584960 458236
rect 583342 458086 584960 458146
rect 583342 458010 583402 458086
rect 583520 458010 584960 458086
rect 583342 457996 584960 458010
rect 583342 457950 583586 457996
rect 61878 456860 61884 456924
rect 61948 456922 61954 456924
rect 583526 456922 583586 457950
rect 61948 456862 583586 456922
rect 61948 456860 61954 456862
rect -960 449578 480 449668
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 2773 423602 2839 423605
rect -960 423600 2839 423602
rect -960 423544 2778 423600
rect 2834 423544 2839 423600
rect -960 423542 2839 423544
rect -960 423452 480 423542
rect 2773 423539 2839 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 582557 365122 582623 365125
rect 583520 365122 584960 365212
rect 582557 365120 584960 365122
rect 582557 365064 582562 365120
rect 582618 365064 584960 365120
rect 582557 365062 584960 365064
rect 582557 365059 582623 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580257 325274 580323 325277
rect 583520 325274 584960 325364
rect 580257 325272 584960 325274
rect 580257 325216 580262 325272
rect 580318 325216 584960 325272
rect 580257 325214 584960 325216
rect 580257 325211 580323 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 68870 313924 68876 313988
rect 68940 313986 68946 313988
rect 75177 313986 75243 313989
rect 68940 313984 75243 313986
rect 68940 313928 75182 313984
rect 75238 313928 75243 313984
rect 68940 313926 75243 313928
rect 68940 313924 68946 313926
rect 75177 313923 75243 313926
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3233 306234 3299 306237
rect -960 306232 3299 306234
rect -960 306176 3238 306232
rect 3294 306176 3299 306232
rect -960 306174 3299 306176
rect -960 306084 480 306174
rect 3233 306171 3299 306174
rect 68645 300930 68711 300933
rect 331254 300930 331260 300932
rect 68645 300928 331260 300930
rect 68645 300872 68650 300928
rect 68706 300872 331260 300928
rect 68645 300870 331260 300872
rect 68645 300867 68711 300870
rect 331254 300868 331260 300870
rect 331324 300868 331330 300932
rect 582649 298754 582715 298757
rect 583520 298754 584960 298844
rect 582649 298752 584960 298754
rect 582649 298696 582654 298752
rect 582710 298696 584960 298752
rect 582649 298694 584960 298696
rect 582649 298691 582715 298694
rect 583520 298604 584960 298694
rect 106089 298210 106155 298213
rect 582465 298210 582531 298213
rect 106089 298208 582531 298210
rect 106089 298152 106094 298208
rect 106150 298152 582470 298208
rect 582526 298152 582531 298208
rect 106089 298150 582531 298152
rect 106089 298147 106155 298150
rect 582465 298147 582531 298150
rect 68829 296850 68895 296853
rect 254526 296850 254532 296852
rect 68829 296848 254532 296850
rect 68829 296792 68834 296848
rect 68890 296792 254532 296848
rect 68829 296790 254532 296792
rect 68829 296787 68895 296790
rect 254526 296788 254532 296790
rect 254596 296788 254602 296852
rect 111793 295490 111859 295493
rect 339493 295490 339559 295493
rect 111793 295488 339559 295490
rect 111793 295432 111798 295488
rect 111854 295432 339498 295488
rect 339554 295432 339559 295488
rect 111793 295430 339559 295432
rect 111793 295427 111859 295430
rect 339493 295427 339559 295430
rect 109953 295354 110019 295357
rect 582925 295354 582991 295357
rect 109953 295352 582991 295354
rect 109953 295296 109958 295352
rect 110014 295296 582930 295352
rect 582986 295296 582991 295352
rect 109953 295294 582991 295296
rect 109953 295291 110019 295294
rect 582925 295291 582991 295294
rect 75821 294266 75887 294269
rect 177297 294266 177363 294269
rect 75821 294264 177363 294266
rect 75821 294208 75826 294264
rect 75882 294208 177302 294264
rect 177358 294208 177363 294264
rect 75821 294206 177363 294208
rect 75821 294203 75887 294206
rect 177297 294203 177363 294206
rect 95785 294130 95851 294133
rect 188337 294130 188403 294133
rect 95785 294128 188403 294130
rect 95785 294072 95790 294128
rect 95846 294072 188342 294128
rect 188398 294072 188403 294128
rect 95785 294070 188403 294072
rect 95785 294067 95851 294070
rect 188337 294067 188403 294070
rect 113173 293994 113239 293997
rect 120022 293994 120028 293996
rect 113173 293992 120028 293994
rect 113173 293936 113178 293992
rect 113234 293936 120028 293992
rect 113173 293934 120028 293936
rect 113173 293931 113239 293934
rect 120022 293932 120028 293934
rect 120092 293932 120098 293996
rect -960 293178 480 293268
rect 2773 293178 2839 293181
rect -960 293176 2839 293178
rect -960 293120 2778 293176
rect 2834 293120 2839 293176
rect -960 293118 2839 293120
rect -960 293028 480 293118
rect 2773 293115 2839 293118
rect 105445 292770 105511 292773
rect 127709 292770 127775 292773
rect 105445 292768 127775 292770
rect 105445 292712 105450 292768
rect 105506 292712 127714 292768
rect 127770 292712 127775 292768
rect 105445 292710 127775 292712
rect 105445 292707 105511 292710
rect 127709 292707 127775 292710
rect 104157 292634 104223 292637
rect 322933 292634 322999 292637
rect 104157 292632 322999 292634
rect 104157 292576 104162 292632
rect 104218 292576 322938 292632
rect 322994 292576 322999 292632
rect 104157 292574 322999 292576
rect 104157 292571 104223 292574
rect 322933 292571 322999 292574
rect 108205 291954 108271 291957
rect 335118 291954 335124 291956
rect 108205 291952 335124 291954
rect 108205 291896 108210 291952
rect 108266 291896 335124 291952
rect 108205 291894 335124 291896
rect 108205 291891 108271 291894
rect 335118 291892 335124 291894
rect 335188 291892 335194 291956
rect 121545 291818 121611 291821
rect 119876 291816 121611 291818
rect 69749 291274 69815 291277
rect 70166 291274 70226 291788
rect 119876 291760 121550 291816
rect 121606 291760 121611 291816
rect 119876 291758 121611 291760
rect 121545 291755 121611 291758
rect 69749 291272 70226 291274
rect 69749 291216 69754 291272
rect 69810 291216 70226 291272
rect 69749 291214 70226 291216
rect 340873 291274 340939 291277
rect 342110 291274 342116 291276
rect 340873 291272 342116 291274
rect 340873 291216 340878 291272
rect 340934 291216 342116 291272
rect 340873 291214 342116 291216
rect 69749 291211 69815 291214
rect 340873 291211 340939 291214
rect 342110 291212 342116 291214
rect 342180 291212 342186 291276
rect 121729 291138 121795 291141
rect 119876 291136 121795 291138
rect 67633 290594 67699 290597
rect 70166 290594 70226 291108
rect 119876 291080 121734 291136
rect 121790 291080 121795 291136
rect 119876 291078 121795 291080
rect 121729 291075 121795 291078
rect 67633 290592 70226 290594
rect 67633 290536 67638 290592
rect 67694 290536 70226 290592
rect 67633 290534 70226 290536
rect 119797 290594 119863 290597
rect 325693 290594 325759 290597
rect 119797 290592 325759 290594
rect 119797 290536 119802 290592
rect 119858 290536 325698 290592
rect 325754 290536 325759 290592
rect 119797 290534 325759 290536
rect 67633 290531 67699 290534
rect 119797 290531 119863 290534
rect 325693 290531 325759 290534
rect 121545 290458 121611 290461
rect 119876 290456 121611 290458
rect 68737 290186 68803 290189
rect 70350 290186 70410 290428
rect 119876 290400 121550 290456
rect 121606 290400 121611 290456
rect 119876 290398 121611 290400
rect 121545 290395 121611 290398
rect 68737 290184 70410 290186
rect 68737 290128 68742 290184
rect 68798 290128 70410 290184
rect 68737 290126 70410 290128
rect 68737 290123 68803 290126
rect 69982 289854 70226 289914
rect 68645 289778 68711 289781
rect 69982 289778 70042 289854
rect 68645 289776 70042 289778
rect 68645 289720 68650 289776
rect 68706 289720 70042 289776
rect 70166 289748 70226 289854
rect 121545 289778 121611 289781
rect 119876 289776 121611 289778
rect 68645 289718 70042 289720
rect 119876 289720 121550 289776
rect 121606 289720 121611 289776
rect 119876 289718 121611 289720
rect 68645 289715 68711 289718
rect 121545 289715 121611 289718
rect 68921 289506 68987 289509
rect 68921 289504 70226 289506
rect 68921 289448 68926 289504
rect 68982 289448 70226 289504
rect 68921 289446 70226 289448
rect 68921 289443 68987 289446
rect 70166 289068 70226 289446
rect 120022 289172 120028 289236
rect 120092 289234 120098 289236
rect 580257 289234 580323 289237
rect 120092 289232 580323 289234
rect 120092 289176 580262 289232
rect 580318 289176 580323 289232
rect 120092 289174 580323 289176
rect 120092 289172 120098 289174
rect 580257 289171 580323 289174
rect 122005 289098 122071 289101
rect 119876 289096 122071 289098
rect 119876 289040 122010 289096
rect 122066 289040 122071 289096
rect 119876 289038 122071 289040
rect 122005 289035 122071 289038
rect 68737 288826 68803 288829
rect 70526 288826 70532 288828
rect 68737 288824 70532 288826
rect 68737 288768 68742 288824
rect 68798 288768 70532 288824
rect 68737 288766 70532 288768
rect 68737 288763 68803 288766
rect 70526 288764 70532 288766
rect 70596 288764 70602 288828
rect 69982 288494 70226 288554
rect 68870 288356 68876 288420
rect 68940 288418 68946 288420
rect 69982 288418 70042 288494
rect 68940 288358 70042 288418
rect 70166 288388 70226 288494
rect 121545 288418 121611 288421
rect 119876 288416 121611 288418
rect 119876 288360 121550 288416
rect 121606 288360 121611 288416
rect 119876 288358 121611 288360
rect 68940 288356 68946 288358
rect 121545 288355 121611 288358
rect 68829 288146 68895 288149
rect 68829 288144 70226 288146
rect 68829 288088 68834 288144
rect 68890 288088 70226 288144
rect 68829 288086 70226 288088
rect 68829 288083 68895 288086
rect 70166 287708 70226 288086
rect 122046 287738 122052 287740
rect 119876 287678 122052 287738
rect 122046 287676 122052 287678
rect 122116 287676 122122 287740
rect 67725 287058 67791 287061
rect 69982 287058 70226 287070
rect 122097 287058 122163 287061
rect 67725 287056 70226 287058
rect 67725 287000 67730 287056
rect 67786 287010 70226 287056
rect 119876 287056 122163 287058
rect 67786 287000 70042 287010
rect 67725 286998 70042 287000
rect 119876 287000 122102 287056
rect 122158 287000 122163 287056
rect 119876 286998 122163 287000
rect 67725 286995 67791 286998
rect 122097 286995 122163 286998
rect 67633 286786 67699 286789
rect 67633 286784 70226 286786
rect 67633 286728 67638 286784
rect 67694 286728 70226 286784
rect 67633 286726 70226 286728
rect 67633 286723 67699 286726
rect 70166 286348 70226 286726
rect 121637 286378 121703 286381
rect 119876 286376 121703 286378
rect 119876 286320 121642 286376
rect 121698 286320 121703 286376
rect 119876 286318 121703 286320
rect 121637 286315 121703 286318
rect 68277 285834 68343 285837
rect 68277 285832 70226 285834
rect 68277 285776 68282 285832
rect 68338 285776 70226 285832
rect 68277 285774 70226 285776
rect 68277 285771 68343 285774
rect 70166 285668 70226 285774
rect 122281 285698 122347 285701
rect 119876 285696 122347 285698
rect 119876 285640 122286 285696
rect 122342 285640 122347 285696
rect 119876 285638 122347 285640
rect 122281 285635 122347 285638
rect 583520 285276 584960 285516
rect 64830 285094 70226 285154
rect 64638 284412 64644 284476
rect 64708 284474 64714 284476
rect 64830 284474 64890 285094
rect 70166 284988 70226 285094
rect 121545 285018 121611 285021
rect 119876 285016 121611 285018
rect 119876 284960 121550 285016
rect 121606 284960 121611 285016
rect 119876 284958 121611 284960
rect 121545 284955 121611 284958
rect 67633 284746 67699 284749
rect 67633 284744 70410 284746
rect 67633 284688 67638 284744
rect 67694 284688 70410 284744
rect 67633 284686 70410 284688
rect 67633 284683 67699 284686
rect 64708 284414 64890 284474
rect 64708 284412 64714 284414
rect 70350 284308 70410 284686
rect 121637 284338 121703 284341
rect 119876 284336 121703 284338
rect 119876 284280 121642 284336
rect 121698 284280 121703 284336
rect 119876 284278 121703 284280
rect 121637 284275 121703 284278
rect 121637 283658 121703 283661
rect 119876 283656 121703 283658
rect 67633 283250 67699 283253
rect 70166 283250 70226 283628
rect 119876 283600 121642 283656
rect 121698 283600 121703 283656
rect 119876 283598 121703 283600
rect 121637 283595 121703 283598
rect 67633 283248 70226 283250
rect 67633 283192 67638 283248
rect 67694 283192 70226 283248
rect 67633 283190 70226 283192
rect 67633 283187 67699 283190
rect 67541 283114 67607 283117
rect 67541 283112 70226 283114
rect 67541 283056 67546 283112
rect 67602 283056 70226 283112
rect 67541 283054 70226 283056
rect 67541 283051 67607 283054
rect 70166 282948 70226 283054
rect 121453 282978 121519 282981
rect 119876 282976 121519 282978
rect 119876 282920 121458 282976
rect 121514 282920 121519 282976
rect 119876 282918 121519 282920
rect 121453 282915 121519 282918
rect 121637 282298 121703 282301
rect 119876 282296 121703 282298
rect 119876 282240 121642 282296
rect 121698 282240 121703 282296
rect 119876 282238 121703 282240
rect 121637 282235 121703 282238
rect 68737 282162 68803 282165
rect 68737 282160 70226 282162
rect 68737 282104 68742 282160
rect 68798 282104 70226 282160
rect 68737 282102 70226 282104
rect 68737 282099 68803 282102
rect 70166 281588 70226 282102
rect 121453 281618 121519 281621
rect 119876 281616 121519 281618
rect 119876 281560 121458 281616
rect 121514 281560 121519 281616
rect 119876 281558 121519 281560
rect 121453 281555 121519 281558
rect 121637 280938 121703 280941
rect 119876 280936 121703 280938
rect 67357 280530 67423 280533
rect 70166 280530 70226 280908
rect 119876 280880 121642 280936
rect 121698 280880 121703 280936
rect 119876 280878 121703 280880
rect 121637 280875 121703 280878
rect 67357 280528 70226 280530
rect 67357 280472 67362 280528
rect 67418 280472 70226 280528
rect 67357 280470 70226 280472
rect 67357 280467 67423 280470
rect 67633 280394 67699 280397
rect 67633 280392 70226 280394
rect 67633 280336 67638 280392
rect 67694 280336 70226 280392
rect 67633 280334 70226 280336
rect 67633 280331 67699 280334
rect 70166 280228 70226 280334
rect 121453 280258 121519 280261
rect 119876 280256 121519 280258
rect -960 279972 480 280212
rect 119876 280200 121458 280256
rect 121514 280200 121519 280256
rect 119876 280198 121519 280200
rect 121453 280195 121519 280198
rect 121637 279578 121703 279581
rect 119876 279576 121703 279578
rect 67633 279170 67699 279173
rect 70166 279170 70226 279548
rect 119876 279520 121642 279576
rect 121698 279520 121703 279576
rect 119876 279518 121703 279520
rect 121637 279515 121703 279518
rect 67633 279168 70226 279170
rect 67633 279112 67638 279168
rect 67694 279112 70226 279168
rect 67633 279110 70226 279112
rect 67633 279107 67699 279110
rect 67725 279034 67791 279037
rect 67725 279032 70226 279034
rect 67725 278976 67730 279032
rect 67786 278976 70226 279032
rect 67725 278974 70226 278976
rect 67725 278971 67791 278974
rect 70166 278868 70226 278974
rect 121453 278898 121519 278901
rect 119876 278896 121519 278898
rect 119876 278840 121458 278896
rect 121514 278840 121519 278896
rect 119876 278838 121519 278840
rect 121453 278835 121519 278838
rect 121637 278218 121703 278221
rect 119876 278216 121703 278218
rect 67725 277810 67791 277813
rect 70166 277810 70226 278188
rect 119876 278160 121642 278216
rect 121698 278160 121703 278216
rect 119876 278158 121703 278160
rect 121637 278155 121703 278158
rect 67725 277808 70226 277810
rect 67725 277752 67730 277808
rect 67786 277752 70226 277808
rect 67725 277750 70226 277752
rect 67725 277747 67791 277750
rect 67633 277674 67699 277677
rect 67633 277672 70226 277674
rect 67633 277616 67638 277672
rect 67694 277616 70226 277672
rect 67633 277614 70226 277616
rect 67633 277611 67699 277614
rect 70166 277508 70226 277614
rect 121453 277538 121519 277541
rect 119876 277536 121519 277538
rect 119876 277480 121458 277536
rect 121514 277480 121519 277536
rect 119876 277478 121519 277480
rect 121453 277475 121519 277478
rect 121453 276858 121519 276861
rect 119876 276856 121519 276858
rect 67633 276450 67699 276453
rect 70166 276450 70226 276828
rect 119876 276800 121458 276856
rect 121514 276800 121519 276856
rect 119876 276798 121519 276800
rect 121453 276795 121519 276798
rect 67633 276448 70226 276450
rect 67633 276392 67638 276448
rect 67694 276392 70226 276448
rect 67633 276390 70226 276392
rect 67633 276387 67699 276390
rect 68001 276314 68067 276317
rect 68001 276312 70226 276314
rect 68001 276256 68006 276312
rect 68062 276256 70226 276312
rect 68001 276254 70226 276256
rect 68001 276251 68067 276254
rect 70166 276148 70226 276254
rect 121637 276178 121703 276181
rect 119876 276176 121703 276178
rect 119876 276120 121642 276176
rect 121698 276120 121703 276176
rect 119876 276118 121703 276120
rect 121637 276115 121703 276118
rect 122097 275498 122163 275501
rect 119876 275496 122163 275498
rect 68369 275226 68435 275229
rect 70166 275226 70226 275468
rect 119876 275440 122102 275496
rect 122158 275440 122163 275496
rect 119876 275438 122163 275440
rect 122097 275435 122163 275438
rect 68369 275224 70226 275226
rect 68369 275168 68374 275224
rect 68430 275168 70226 275224
rect 68369 275166 70226 275168
rect 68369 275163 68435 275166
rect 67633 275090 67699 275093
rect 67633 275088 70410 275090
rect 67633 275032 67638 275088
rect 67694 275032 70410 275088
rect 67633 275030 70410 275032
rect 67633 275027 67699 275030
rect 70350 274788 70410 275030
rect 121453 274818 121519 274821
rect 119876 274816 121519 274818
rect 119876 274760 121458 274816
rect 121514 274760 121519 274816
rect 119876 274758 121519 274760
rect 121453 274755 121519 274758
rect 67725 274546 67791 274549
rect 67725 274544 70226 274546
rect 67725 274488 67730 274544
rect 67786 274488 70226 274544
rect 67725 274486 70226 274488
rect 67725 274483 67791 274486
rect 70166 274108 70226 274486
rect 121453 274138 121519 274141
rect 119876 274136 121519 274138
rect 119876 274080 121458 274136
rect 121514 274080 121519 274136
rect 119876 274078 121519 274080
rect 121453 274075 121519 274078
rect 68001 273594 68067 273597
rect 68001 273592 70226 273594
rect 68001 273536 68006 273592
rect 68062 273536 70226 273592
rect 68001 273534 70226 273536
rect 68001 273531 68067 273534
rect 70166 273428 70226 273534
rect 121453 273458 121519 273461
rect 119876 273456 121519 273458
rect 119876 273400 121458 273456
rect 121514 273400 121519 273456
rect 119876 273398 121519 273400
rect 121453 273395 121519 273398
rect 121545 272778 121611 272781
rect 119876 272776 121611 272778
rect 67725 272370 67791 272373
rect 70166 272370 70226 272748
rect 119876 272720 121550 272776
rect 121606 272720 121611 272776
rect 119876 272718 121611 272720
rect 121545 272715 121611 272718
rect 67725 272368 70226 272370
rect 67725 272312 67730 272368
rect 67786 272312 70226 272368
rect 67725 272310 70226 272312
rect 67725 272307 67791 272310
rect 67633 272234 67699 272237
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 67633 272232 70226 272234
rect 67633 272176 67638 272232
rect 67694 272176 70226 272232
rect 67633 272174 70226 272176
rect 67633 272171 67699 272174
rect 70166 272068 70226 272174
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 119876 272038 122850 272098
rect 583520 272084 584960 272174
rect 122790 271962 122850 272038
rect 166942 271962 166948 271964
rect 122790 271902 166948 271962
rect 166942 271900 166948 271902
rect 167012 271900 167018 271964
rect 121545 271418 121611 271421
rect 119876 271416 121611 271418
rect 67633 271010 67699 271013
rect 70166 271010 70226 271388
rect 119876 271360 121550 271416
rect 121606 271360 121611 271416
rect 119876 271358 121611 271360
rect 121545 271355 121611 271358
rect 67633 271008 70226 271010
rect 67633 270952 67638 271008
rect 67694 270952 70226 271008
rect 67633 270950 70226 270952
rect 67633 270947 67699 270950
rect 69013 270874 69079 270877
rect 69013 270872 70226 270874
rect 69013 270816 69018 270872
rect 69074 270816 70226 270872
rect 69013 270814 70226 270816
rect 69013 270811 69079 270814
rect 70166 270708 70226 270814
rect 121453 270058 121519 270061
rect 119876 270056 121519 270058
rect 67633 269650 67699 269653
rect 70166 269650 70226 270028
rect 119876 270000 121458 270056
rect 121514 270000 121519 270056
rect 119876 269998 121519 270000
rect 121453 269995 121519 269998
rect 122046 269724 122052 269788
rect 122116 269786 122122 269788
rect 392577 269786 392643 269789
rect 122116 269784 392643 269786
rect 122116 269728 392582 269784
rect 392638 269728 392643 269784
rect 122116 269726 392643 269728
rect 122116 269724 122122 269726
rect 392577 269723 392643 269726
rect 67633 269648 70226 269650
rect 67633 269592 67638 269648
rect 67694 269592 70226 269648
rect 67633 269590 70226 269592
rect 67633 269587 67699 269590
rect 67265 269514 67331 269517
rect 67265 269512 70226 269514
rect 67265 269456 67270 269512
rect 67326 269456 70226 269512
rect 67265 269454 70226 269456
rect 67265 269451 67331 269454
rect 70166 269348 70226 269454
rect 119876 269318 122850 269378
rect 122790 269242 122850 269318
rect 263542 269242 263548 269244
rect 122790 269182 263548 269242
rect 263542 269180 263548 269182
rect 263612 269180 263618 269244
rect 120073 268698 120139 268701
rect 119876 268696 120139 268698
rect 69197 268290 69263 268293
rect 70166 268290 70226 268668
rect 119876 268640 120078 268696
rect 120134 268640 120139 268696
rect 119876 268638 120139 268640
rect 120073 268635 120139 268638
rect 69197 268288 70226 268290
rect 69197 268232 69202 268288
rect 69258 268232 70226 268288
rect 69197 268230 70226 268232
rect 69197 268227 69263 268230
rect 67633 268154 67699 268157
rect 67633 268152 70226 268154
rect 67633 268096 67638 268152
rect 67694 268096 70226 268152
rect 67633 268094 70226 268096
rect 67633 268091 67699 268094
rect 70166 267988 70226 268094
rect 121453 268018 121519 268021
rect 119876 268016 121519 268018
rect 119876 267960 121458 268016
rect 121514 267960 121519 268016
rect 119876 267958 121519 267960
rect 121453 267955 121519 267958
rect 67725 267474 67791 267477
rect 67725 267472 70226 267474
rect 67725 267416 67730 267472
rect 67786 267416 70226 267472
rect 67725 267414 70226 267416
rect 67725 267411 67791 267414
rect 70166 267308 70226 267414
rect 121545 267338 121611 267341
rect 119876 267336 121611 267338
rect -960 267202 480 267292
rect 119876 267280 121550 267336
rect 121606 267280 121611 267336
rect 119876 267278 121611 267280
rect 121545 267275 121611 267278
rect 3601 267202 3667 267205
rect -960 267200 3667 267202
rect -960 267144 3606 267200
rect 3662 267144 3667 267200
rect -960 267142 3667 267144
rect -960 267052 480 267142
rect 3601 267139 3667 267142
rect 67633 267066 67699 267069
rect 67633 267064 70226 267066
rect 67633 267008 67638 267064
rect 67694 267008 70226 267064
rect 67633 267006 70226 267008
rect 67633 267003 67699 267006
rect 70166 266628 70226 267006
rect 121453 266658 121519 266661
rect 119876 266656 121519 266658
rect 119876 266600 121458 266656
rect 121514 266600 121519 266656
rect 119876 266598 121519 266600
rect 121453 266595 121519 266598
rect 121545 265978 121611 265981
rect 119876 265976 121611 265978
rect 67633 265434 67699 265437
rect 70166 265434 70226 265948
rect 119876 265920 121550 265976
rect 121606 265920 121611 265976
rect 119876 265918 121611 265920
rect 121545 265915 121611 265918
rect 67633 265432 70226 265434
rect 67633 265376 67638 265432
rect 67694 265376 70226 265432
rect 67633 265374 70226 265376
rect 67633 265371 67699 265374
rect 121453 265298 121519 265301
rect 119876 265296 121519 265298
rect 67725 265026 67791 265029
rect 70350 265026 70410 265268
rect 119876 265240 121458 265296
rect 121514 265240 121519 265296
rect 119876 265238 121519 265240
rect 121453 265235 121519 265238
rect 67725 265024 70410 265026
rect 67725 264968 67730 265024
rect 67786 264968 70410 265024
rect 67725 264966 70410 264968
rect 67725 264963 67791 264966
rect 121637 264618 121703 264621
rect 119876 264616 121703 264618
rect 67725 264210 67791 264213
rect 70166 264210 70226 264588
rect 119876 264560 121642 264616
rect 121698 264560 121703 264616
rect 119876 264558 121703 264560
rect 121637 264555 121703 264558
rect 67725 264208 70226 264210
rect 67725 264152 67730 264208
rect 67786 264152 70226 264208
rect 67725 264150 70226 264152
rect 122097 264210 122163 264213
rect 340086 264210 340092 264212
rect 122097 264208 340092 264210
rect 122097 264152 122102 264208
rect 122158 264152 340092 264208
rect 122097 264150 340092 264152
rect 67725 264147 67791 264150
rect 122097 264147 122163 264150
rect 340086 264148 340092 264150
rect 340156 264148 340162 264212
rect 121545 263938 121611 263941
rect 119876 263936 121611 263938
rect 67633 263666 67699 263669
rect 70350 263666 70410 263908
rect 119876 263880 121550 263936
rect 121606 263880 121611 263936
rect 119876 263878 121611 263880
rect 121545 263875 121611 263878
rect 67633 263664 70410 263666
rect 67633 263608 67638 263664
rect 67694 263608 70410 263664
rect 67633 263606 70410 263608
rect 67633 263603 67699 263606
rect 67633 263530 67699 263533
rect 67633 263528 70226 263530
rect 67633 263472 67638 263528
rect 67694 263472 70226 263528
rect 67633 263470 70226 263472
rect 67633 263467 67699 263470
rect 70166 263228 70226 263470
rect 121453 263258 121519 263261
rect 119876 263256 121519 263258
rect 119876 263200 121458 263256
rect 121514 263200 121519 263256
rect 119876 263198 121519 263200
rect 121453 263195 121519 263198
rect 121453 262578 121519 262581
rect 119876 262576 121519 262578
rect 67633 262306 67699 262309
rect 70166 262306 70226 262548
rect 119876 262520 121458 262576
rect 121514 262520 121519 262576
rect 119876 262518 121519 262520
rect 121453 262515 121519 262518
rect 67633 262304 70226 262306
rect 67633 262248 67638 262304
rect 67694 262248 70226 262304
rect 67633 262246 70226 262248
rect 67633 262243 67699 262246
rect 121453 261898 121519 261901
rect 119876 261896 121519 261898
rect 67725 261490 67791 261493
rect 70166 261490 70226 261868
rect 119876 261840 121458 261896
rect 121514 261840 121519 261896
rect 119876 261838 121519 261840
rect 121453 261835 121519 261838
rect 67725 261488 70226 261490
rect 67725 261432 67730 261488
rect 67786 261432 70226 261488
rect 67725 261430 70226 261432
rect 67725 261427 67791 261430
rect 120257 261218 120323 261221
rect 119876 261216 120323 261218
rect 67633 260946 67699 260949
rect 70350 260946 70410 261188
rect 119876 261160 120262 261216
rect 120318 261160 120323 261216
rect 119876 261158 120323 261160
rect 120257 261155 120323 261158
rect 67633 260944 70410 260946
rect 67633 260888 67638 260944
rect 67694 260888 70410 260944
rect 67633 260886 70410 260888
rect 67633 260883 67699 260886
rect 67633 260810 67699 260813
rect 67633 260808 70226 260810
rect 67633 260752 67638 260808
rect 67694 260752 70226 260808
rect 67633 260750 70226 260752
rect 67633 260747 67699 260750
rect 70166 260508 70226 260750
rect 119846 259994 119906 260508
rect 119846 259934 122850 259994
rect 121453 259858 121519 259861
rect 119876 259856 121519 259858
rect 67633 259586 67699 259589
rect 70350 259586 70410 259828
rect 119876 259800 121458 259856
rect 121514 259800 121519 259856
rect 119876 259798 121519 259800
rect 121453 259795 121519 259798
rect 67633 259584 70410 259586
rect 67633 259528 67638 259584
rect 67694 259528 70410 259584
rect 67633 259526 70410 259528
rect 122790 259586 122850 259934
rect 338614 259586 338620 259588
rect 122790 259526 338620 259586
rect 67633 259523 67699 259526
rect 338614 259524 338620 259526
rect 338684 259524 338690 259588
rect 121453 259178 121519 259181
rect 119876 259176 121519 259178
rect 67725 258634 67791 258637
rect 70166 258634 70226 259148
rect 119876 259120 121458 259176
rect 121514 259120 121519 259176
rect 119876 259118 121519 259120
rect 121453 259115 121519 259118
rect 579797 258906 579863 258909
rect 583520 258906 584960 258996
rect 579797 258904 584960 258906
rect 579797 258848 579802 258904
rect 579858 258848 584960 258904
rect 579797 258846 584960 258848
rect 579797 258843 579863 258846
rect 583520 258756 584960 258846
rect 67725 258632 70226 258634
rect 67725 258576 67730 258632
rect 67786 258576 70226 258632
rect 67725 258574 70226 258576
rect 67725 258571 67791 258574
rect 121545 258498 121611 258501
rect 119876 258496 121611 258498
rect 67633 258226 67699 258229
rect 70166 258226 70226 258468
rect 119876 258440 121550 258496
rect 121606 258440 121611 258496
rect 119876 258438 121611 258440
rect 121545 258435 121611 258438
rect 67633 258224 70226 258226
rect 67633 258168 67638 258224
rect 67694 258168 70226 258224
rect 67633 258166 70226 258168
rect 67633 258163 67699 258166
rect 121545 257818 121611 257821
rect 119876 257816 121611 257818
rect 67633 257274 67699 257277
rect 70166 257274 70226 257788
rect 119876 257760 121550 257816
rect 121606 257760 121611 257816
rect 119876 257758 121611 257760
rect 121545 257755 121611 257758
rect 67633 257272 70226 257274
rect 67633 257216 67638 257272
rect 67694 257216 70226 257272
rect 67633 257214 70226 257216
rect 67633 257211 67699 257214
rect 121453 257138 121519 257141
rect 119876 257136 121519 257138
rect 66110 256668 66116 256732
rect 66180 256730 66186 256732
rect 70166 256730 70226 257108
rect 119876 257080 121458 257136
rect 121514 257080 121519 257136
rect 119876 257078 121519 257080
rect 121453 257075 121519 257078
rect 66180 256670 70226 256730
rect 66180 256668 66186 256670
rect 121453 256458 121519 256461
rect 119876 256456 121519 256458
rect 67633 255914 67699 255917
rect 70166 255914 70226 256428
rect 119876 256400 121458 256456
rect 121514 256400 121519 256456
rect 119876 256398 121519 256400
rect 121453 256395 121519 256398
rect 67633 255912 70226 255914
rect 67633 255856 67638 255912
rect 67694 255856 70226 255912
rect 67633 255854 70226 255856
rect 67633 255851 67699 255854
rect 121637 255778 121703 255781
rect 119876 255776 121703 255778
rect 67725 255370 67791 255373
rect 70166 255370 70226 255748
rect 119876 255720 121642 255776
rect 121698 255720 121703 255776
rect 119876 255718 121703 255720
rect 121637 255715 121703 255718
rect 67725 255368 70226 255370
rect 67725 255312 67730 255368
rect 67786 255312 70226 255368
rect 67725 255310 70226 255312
rect 67725 255307 67791 255310
rect 67633 255234 67699 255237
rect 67633 255232 70226 255234
rect 67633 255176 67638 255232
rect 67694 255176 70226 255232
rect 67633 255174 70226 255176
rect 67633 255171 67699 255174
rect 70166 255068 70226 255174
rect 121545 255098 121611 255101
rect 119876 255096 121611 255098
rect 119876 255040 121550 255096
rect 121606 255040 121611 255096
rect 119876 255038 121611 255040
rect 121545 255035 121611 255038
rect 121453 254418 121519 254421
rect 119876 254416 121519 254418
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 62982 254084 62988 254148
rect 63052 254146 63058 254148
rect 70166 254146 70226 254388
rect 119876 254360 121458 254416
rect 121514 254360 121519 254416
rect 119876 254358 121519 254360
rect 121453 254355 121519 254358
rect 63052 254086 70226 254146
rect 63052 254084 63058 254086
rect 122097 253738 122163 253741
rect 119876 253736 122163 253738
rect 67725 253194 67791 253197
rect 70166 253194 70226 253708
rect 119876 253680 122102 253736
rect 122158 253680 122163 253736
rect 119876 253678 122163 253680
rect 122097 253675 122163 253678
rect 67725 253192 70226 253194
rect 67725 253136 67730 253192
rect 67786 253136 70226 253192
rect 67725 253134 70226 253136
rect 67725 253131 67791 253134
rect 120022 253132 120028 253196
rect 120092 253194 120098 253196
rect 142797 253194 142863 253197
rect 120092 253192 142863 253194
rect 120092 253136 142802 253192
rect 142858 253136 142863 253192
rect 120092 253134 142863 253136
rect 120092 253132 120098 253134
rect 142797 253131 142863 253134
rect 121545 253058 121611 253061
rect 119876 253056 121611 253058
rect 67633 252786 67699 252789
rect 70350 252786 70410 253028
rect 119876 253000 121550 253056
rect 121606 253000 121611 253056
rect 119876 252998 121611 253000
rect 121545 252995 121611 252998
rect 67633 252784 70410 252786
rect 67633 252728 67638 252784
rect 67694 252728 70410 252784
rect 67633 252726 70410 252728
rect 67633 252723 67699 252726
rect 121453 252378 121519 252381
rect 119876 252376 121519 252378
rect 67633 251834 67699 251837
rect 70166 251834 70226 252348
rect 119876 252320 121458 252376
rect 121514 252320 121519 252376
rect 119876 252318 121519 252320
rect 121453 252315 121519 252318
rect 67633 251832 70226 251834
rect 67633 251776 67638 251832
rect 67694 251776 70226 251832
rect 67633 251774 70226 251776
rect 67633 251771 67699 251774
rect 121453 251698 121519 251701
rect 119876 251696 121519 251698
rect 69105 251290 69171 251293
rect 70166 251290 70226 251668
rect 119876 251640 121458 251696
rect 121514 251640 121519 251696
rect 119876 251638 121519 251640
rect 121453 251635 121519 251638
rect 69105 251288 70226 251290
rect 69105 251232 69110 251288
rect 69166 251232 70226 251288
rect 69105 251230 70226 251232
rect 69105 251227 69171 251230
rect 120073 251018 120139 251021
rect 119876 251016 120139 251018
rect 67725 250474 67791 250477
rect 70166 250474 70226 250988
rect 119876 250960 120078 251016
rect 120134 250960 120139 251016
rect 119876 250958 120139 250960
rect 120073 250955 120139 250958
rect 67725 250472 70226 250474
rect 67725 250416 67730 250472
rect 67786 250416 70226 250472
rect 67725 250414 70226 250416
rect 67725 250411 67791 250414
rect 121545 250338 121611 250341
rect 119876 250336 121611 250338
rect 67633 249930 67699 249933
rect 70166 249930 70226 250308
rect 119876 250280 121550 250336
rect 121606 250280 121611 250336
rect 119876 250278 121611 250280
rect 121545 250275 121611 250278
rect 67633 249928 70226 249930
rect 67633 249872 67638 249928
rect 67694 249872 70226 249928
rect 67633 249870 70226 249872
rect 67633 249867 67699 249870
rect 67633 249794 67699 249797
rect 67633 249792 70226 249794
rect 67633 249736 67638 249792
rect 67694 249736 70226 249792
rect 67633 249734 70226 249736
rect 67633 249731 67699 249734
rect 70166 249628 70226 249734
rect 121453 249658 121519 249661
rect 119876 249656 121519 249658
rect 119876 249600 121458 249656
rect 121514 249600 121519 249656
rect 119876 249598 121519 249600
rect 121453 249595 121519 249598
rect 121453 248978 121519 248981
rect 119876 248976 121519 248978
rect 67633 248570 67699 248573
rect 70166 248570 70226 248948
rect 119876 248920 121458 248976
rect 121514 248920 121519 248976
rect 119876 248918 121519 248920
rect 121453 248915 121519 248918
rect 67633 248568 70226 248570
rect 67633 248512 67638 248568
rect 67694 248512 70226 248568
rect 67633 248510 70226 248512
rect 67633 248507 67699 248510
rect 121453 248298 121519 248301
rect 119876 248296 121519 248298
rect 67633 247754 67699 247757
rect 70166 247754 70226 248268
rect 119876 248240 121458 248296
rect 121514 248240 121519 248296
rect 119876 248238 121519 248240
rect 121453 248235 121519 248238
rect 67633 247752 70226 247754
rect 67633 247696 67638 247752
rect 67694 247696 70226 247752
rect 67633 247694 70226 247696
rect 67633 247691 67699 247694
rect 120165 247618 120231 247621
rect 119876 247616 120231 247618
rect 67725 247210 67791 247213
rect 70166 247210 70226 247588
rect 119876 247560 120170 247616
rect 120226 247560 120231 247616
rect 119876 247558 120231 247560
rect 120165 247555 120231 247558
rect 67725 247208 70226 247210
rect 67725 247152 67730 247208
rect 67786 247152 70226 247208
rect 67725 247150 70226 247152
rect 67725 247147 67791 247150
rect 121545 246938 121611 246941
rect 119876 246936 121611 246938
rect 67633 246666 67699 246669
rect 70350 246666 70410 246908
rect 119876 246880 121550 246936
rect 121606 246880 121611 246936
rect 119876 246878 121611 246880
rect 121545 246875 121611 246878
rect 67633 246664 70410 246666
rect 67633 246608 67638 246664
rect 67694 246608 70410 246664
rect 67633 246606 70410 246608
rect 67633 246603 67699 246606
rect 67725 245986 67791 245989
rect 70166 245986 70226 246228
rect 67725 245984 70226 245986
rect 67725 245928 67730 245984
rect 67786 245928 70226 245984
rect 67725 245926 70226 245928
rect 67725 245923 67791 245926
rect 119846 245714 119906 246228
rect 258390 245714 258396 245716
rect 119846 245654 258396 245714
rect 258390 245652 258396 245654
rect 258460 245652 258466 245716
rect 121545 245578 121611 245581
rect 119876 245576 121611 245578
rect 67633 245306 67699 245309
rect 70350 245306 70410 245548
rect 119876 245520 121550 245576
rect 121606 245520 121611 245576
rect 119876 245518 121611 245520
rect 121545 245515 121611 245518
rect 579889 245578 579955 245581
rect 583520 245578 584960 245668
rect 579889 245576 584960 245578
rect 579889 245520 579894 245576
rect 579950 245520 584960 245576
rect 579889 245518 584960 245520
rect 579889 245515 579955 245518
rect 583520 245428 584960 245518
rect 67633 245304 70410 245306
rect 67633 245248 67638 245304
rect 67694 245248 70410 245304
rect 67633 245246 70410 245248
rect 67633 245243 67699 245246
rect 121453 244898 121519 244901
rect 119876 244896 121519 244898
rect 67633 244626 67699 244629
rect 70166 244626 70226 244868
rect 119876 244840 121458 244896
rect 121514 244840 121519 244896
rect 119876 244838 121519 244840
rect 121453 244835 121519 244838
rect 67633 244624 70226 244626
rect 67633 244568 67638 244624
rect 67694 244568 70226 244624
rect 67633 244566 70226 244568
rect 67633 244563 67699 244566
rect 69982 244294 70226 244354
rect 69657 244218 69723 244221
rect 69982 244218 70042 244294
rect 69657 244216 70042 244218
rect 69657 244160 69662 244216
rect 69718 244160 70042 244216
rect 70166 244188 70226 244294
rect 121637 244218 121703 244221
rect 119876 244216 121703 244218
rect 69657 244158 70042 244160
rect 119876 244160 121642 244216
rect 121698 244160 121703 244216
rect 119876 244158 121703 244160
rect 69657 244155 69723 244158
rect 121637 244155 121703 244158
rect 67725 243946 67791 243949
rect 67725 243944 70226 243946
rect 67725 243888 67730 243944
rect 67786 243888 70226 243944
rect 67725 243886 70226 243888
rect 67725 243883 67791 243886
rect 70166 243508 70226 243886
rect 121453 243538 121519 243541
rect 119876 243536 121519 243538
rect 119876 243480 121458 243536
rect 121514 243480 121519 243536
rect 119876 243478 121519 243480
rect 121453 243475 121519 243478
rect 121453 242858 121519 242861
rect 119876 242856 121519 242858
rect 70166 242314 70226 242828
rect 119876 242800 121458 242856
rect 121514 242800 121519 242856
rect 119876 242798 121519 242800
rect 121453 242795 121519 242798
rect 64830 242254 70226 242314
rect 59118 241708 59124 241772
rect 59188 241770 59194 241772
rect 64830 241770 64890 242254
rect 121545 242178 121611 242181
rect 119876 242176 121611 242178
rect 67633 241906 67699 241909
rect 70166 241906 70226 242148
rect 119876 242120 121550 242176
rect 121606 242120 121611 242176
rect 119876 242118 121611 242120
rect 121545 242115 121611 242118
rect 67633 241904 70226 241906
rect 67633 241848 67638 241904
rect 67694 241848 70226 241904
rect 67633 241846 70226 241848
rect 67633 241843 67699 241846
rect 59188 241710 64890 241770
rect 59188 241708 59194 241710
rect -960 241090 480 241180
rect 3049 241090 3115 241093
rect -960 241088 3115 241090
rect -960 241032 3054 241088
rect 3110 241032 3115 241088
rect -960 241030 3115 241032
rect -960 240940 480 241030
rect 3049 241027 3115 241030
rect 70166 240954 70226 241468
rect 119846 240957 119906 241468
rect 64830 240894 70226 240954
rect 119797 240952 119906 240957
rect 119797 240896 119802 240952
rect 119858 240896 119906 240952
rect 119797 240894 119906 240896
rect 61878 240348 61884 240412
rect 61948 240410 61954 240412
rect 64830 240410 64890 240894
rect 119797 240891 119863 240894
rect 121453 240818 121519 240821
rect 119876 240816 121519 240818
rect 61948 240350 64890 240410
rect 61948 240348 61954 240350
rect 67449 240274 67515 240277
rect 70166 240274 70226 240788
rect 119876 240760 121458 240816
rect 121514 240760 121519 240816
rect 119876 240758 121519 240760
rect 121453 240755 121519 240758
rect 67449 240272 70226 240274
rect 67449 240216 67454 240272
rect 67510 240216 70226 240272
rect 67449 240214 70226 240216
rect 67449 240211 67515 240214
rect 121545 240138 121611 240141
rect 119876 240136 121611 240138
rect 119876 240080 121550 240136
rect 121606 240080 121611 240136
rect 119876 240078 121611 240080
rect 121545 240075 121611 240078
rect 118969 239866 119035 239869
rect 120022 239866 120028 239868
rect 118969 239864 120028 239866
rect 118969 239808 118974 239864
rect 119030 239808 120028 239864
rect 118969 239806 120028 239808
rect 118969 239803 119035 239806
rect 120022 239804 120028 239806
rect 120092 239804 120098 239868
rect 66110 236540 66116 236604
rect 66180 236602 66186 236604
rect 345054 236602 345060 236604
rect 66180 236542 345060 236602
rect 66180 236540 66186 236542
rect 345054 236540 345060 236542
rect 345124 236540 345130 236604
rect 62982 232460 62988 232524
rect 63052 232522 63058 232524
rect 582833 232522 582899 232525
rect 63052 232520 582899 232522
rect 63052 232464 582838 232520
rect 582894 232464 582899 232520
rect 63052 232462 582899 232464
rect 63052 232460 63058 232462
rect 582833 232459 582899 232462
rect 580349 232386 580415 232389
rect 583520 232386 584960 232476
rect 580349 232384 584960 232386
rect 580349 232328 580354 232384
rect 580410 232328 584960 232384
rect 580349 232326 584960 232328
rect 580349 232323 580415 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 64638 226884 64644 226948
rect 64708 226946 64714 226948
rect 574737 226946 574803 226949
rect 64708 226944 574803 226946
rect 64708 226888 574742 226944
rect 574798 226888 574803 226944
rect 64708 226886 574803 226888
rect 64708 226884 64714 226886
rect 574737 226883 574803 226886
rect 73245 225586 73311 225589
rect 320214 225586 320220 225588
rect 73245 225584 320220 225586
rect 73245 225528 73250 225584
rect 73306 225528 320220 225584
rect 73245 225526 320220 225528
rect 73245 225523 73311 225526
rect 320214 225524 320220 225526
rect 320284 225524 320290 225588
rect 84377 222866 84443 222869
rect 327022 222866 327028 222868
rect 84377 222864 327028 222866
rect 84377 222808 84382 222864
rect 84438 222808 327028 222864
rect 84377 222806 327028 222808
rect 84377 222803 84443 222806
rect 327022 222804 327028 222806
rect 327092 222804 327098 222868
rect 583017 219058 583083 219061
rect 583520 219058 584960 219148
rect 583017 219056 584960 219058
rect 583017 219000 583022 219056
rect 583078 219000 584960 219056
rect 583017 218998 584960 219000
rect 583017 218995 583083 218998
rect 583520 218908 584960 218998
rect 59077 218650 59143 218653
rect 267774 218650 267780 218652
rect 59077 218648 267780 218650
rect 59077 218592 59082 218648
rect 59138 218592 267780 218648
rect 59077 218590 267780 218592
rect 59077 218587 59143 218590
rect 267774 218588 267780 218590
rect 267844 218588 267850 218652
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 114553 213210 114619 213213
rect 327206 213210 327212 213212
rect 114553 213208 327212 213210
rect 114553 213152 114558 213208
rect 114614 213152 327212 213208
rect 114553 213150 327212 213152
rect 114553 213147 114619 213150
rect 327206 213148 327212 213150
rect 327276 213148 327282 213212
rect 50981 211850 51047 211853
rect 342294 211850 342300 211852
rect 50981 211848 342300 211850
rect 50981 211792 50986 211848
rect 51042 211792 342300 211848
rect 50981 211790 342300 211792
rect 50981 211787 51047 211790
rect 342294 211788 342300 211790
rect 342364 211788 342370 211852
rect 49601 210354 49667 210357
rect 334014 210354 334020 210356
rect 49601 210352 334020 210354
rect 49601 210296 49606 210352
rect 49662 210296 334020 210352
rect 49601 210294 334020 210296
rect 49601 210291 49667 210294
rect 334014 210292 334020 210294
rect 334084 210292 334090 210356
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect 64597 203554 64663 203557
rect 269062 203554 269068 203556
rect 64597 203552 269068 203554
rect 64597 203496 64602 203552
rect 64658 203496 269068 203552
rect 64597 203494 269068 203496
rect 64597 203491 64663 203494
rect 269062 203492 269068 203494
rect 269132 203492 269138 203556
rect -960 201922 480 202012
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 69105 196618 69171 196621
rect 324262 196618 324268 196620
rect 69105 196616 324268 196618
rect 69105 196560 69110 196616
rect 69166 196560 324268 196616
rect 69105 196558 324268 196560
rect 69105 196555 69171 196558
rect 324262 196556 324268 196558
rect 324332 196556 324338 196620
rect 334617 194578 334683 194581
rect 336774 194578 336780 194580
rect 334617 194576 336780 194578
rect 334617 194520 334622 194576
rect 334678 194520 336780 194576
rect 334617 194518 336780 194520
rect 334617 194515 334683 194518
rect 336774 194516 336780 194518
rect 336844 194516 336850 194580
rect 79317 192538 79383 192541
rect 266302 192538 266308 192540
rect 79317 192536 266308 192538
rect 79317 192480 79322 192536
rect 79378 192480 266308 192536
rect 79317 192478 266308 192480
rect 79317 192475 79383 192478
rect 266302 192476 266308 192478
rect 266372 192476 266378 192540
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect 62021 191042 62087 191045
rect 263726 191042 263732 191044
rect 62021 191040 263732 191042
rect 62021 190984 62026 191040
rect 62082 190984 263732 191040
rect 62021 190982 263732 190984
rect 62021 190979 62087 190982
rect 263726 190980 263732 190982
rect 263796 190980 263802 191044
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 92473 188322 92539 188325
rect 342437 188322 342503 188325
rect 92473 188320 342503 188322
rect 92473 188264 92478 188320
rect 92534 188264 342442 188320
rect 342498 188264 342503 188320
rect 92473 188262 342503 188264
rect 92473 188259 92539 188262
rect 342437 188259 342503 188262
rect 197997 185602 198063 185605
rect 256734 185602 256740 185604
rect 197997 185600 256740 185602
rect 197997 185544 198002 185600
rect 198058 185544 256740 185600
rect 197997 185542 256740 185544
rect 197997 185539 198063 185542
rect 256734 185540 256740 185542
rect 256804 185540 256810 185604
rect 99281 183698 99347 183701
rect 166206 183698 166212 183700
rect 99281 183696 166212 183698
rect 99281 183640 99286 183696
rect 99342 183640 166212 183696
rect 99281 183638 166212 183640
rect 99281 183635 99347 183638
rect 166206 183636 166212 183638
rect 166276 183636 166282 183700
rect 71773 182882 71839 182885
rect 341057 182882 341123 182885
rect 71773 182880 341123 182882
rect 71773 182824 71778 182880
rect 71834 182824 341062 182880
rect 341118 182824 341123 182880
rect 71773 182822 341123 182824
rect 71773 182819 71839 182822
rect 341057 182819 341123 182822
rect 59261 180026 59327 180029
rect 335486 180026 335492 180028
rect 59261 180024 335492 180026
rect 59261 179968 59266 180024
rect 59322 179968 335492 180024
rect 59261 179966 335492 179968
rect 59261 179963 59327 179966
rect 335486 179964 335492 179966
rect 335556 179964 335562 180028
rect 110689 179482 110755 179485
rect 166390 179482 166396 179484
rect 110689 179480 166396 179482
rect 110689 179424 110694 179480
rect 110750 179424 166396 179480
rect 110689 179422 166396 179424
rect 110689 179419 110755 179422
rect 166390 179420 166396 179422
rect 166460 179420 166466 179484
rect 338297 179348 338363 179349
rect 338246 179284 338252 179348
rect 338316 179346 338363 179348
rect 338316 179344 338408 179346
rect 338358 179288 338408 179344
rect 338316 179286 338408 179288
rect 338316 179284 338363 179286
rect 338297 179283 338363 179284
rect 582925 179210 582991 179213
rect 583520 179210 584960 179300
rect 582925 179208 584960 179210
rect 582925 179152 582930 179208
rect 582986 179152 584960 179208
rect 582925 179150 584960 179152
rect 582925 179147 582991 179150
rect 583520 179060 584960 179150
rect 302877 178938 302943 178941
rect 334198 178938 334204 178940
rect 302877 178936 334204 178938
rect 302877 178880 302882 178936
rect 302938 178880 334204 178936
rect 302877 178878 334204 178880
rect 302877 178875 302943 178878
rect 334198 178876 334204 178878
rect 334268 178876 334274 178940
rect 245009 178802 245075 178805
rect 255262 178802 255268 178804
rect 245009 178800 255268 178802
rect 245009 178744 245014 178800
rect 245070 178744 255268 178800
rect 245009 178742 255268 178744
rect 245009 178739 245075 178742
rect 255262 178740 255268 178742
rect 255332 178740 255338 178804
rect 298737 178802 298803 178805
rect 332542 178802 332548 178804
rect 298737 178800 332548 178802
rect 298737 178744 298742 178800
rect 298798 178744 332548 178800
rect 298737 178742 332548 178744
rect 298737 178739 298803 178742
rect 332542 178740 332548 178742
rect 332612 178740 332618 178804
rect 60641 178666 60707 178669
rect 328729 178666 328795 178669
rect 60641 178664 328795 178666
rect 60641 178608 60646 178664
rect 60702 178608 328734 178664
rect 328790 178608 328795 178664
rect 60641 178606 328795 178608
rect 60641 178603 60707 178606
rect 328729 178603 328795 178606
rect 97022 177652 97028 177716
rect 97092 177714 97098 177716
rect 97533 177714 97599 177717
rect 97092 177712 97599 177714
rect 97092 177656 97538 177712
rect 97594 177656 97599 177712
rect 97092 177654 97599 177656
rect 97092 177652 97098 177654
rect 97533 177651 97599 177654
rect 98310 177652 98316 177716
rect 98380 177714 98386 177716
rect 99281 177714 99347 177717
rect 98380 177712 99347 177714
rect 98380 177656 99286 177712
rect 99342 177656 99347 177712
rect 98380 177654 99347 177656
rect 98380 177652 98386 177654
rect 99281 177651 99347 177654
rect 105670 177652 105676 177716
rect 105740 177714 105746 177716
rect 106181 177714 106247 177717
rect 105740 177712 106247 177714
rect 105740 177656 106186 177712
rect 106242 177656 106247 177712
rect 105740 177654 106247 177656
rect 105740 177652 105746 177654
rect 106181 177651 106247 177654
rect 106958 177652 106964 177716
rect 107028 177714 107034 177716
rect 107561 177714 107627 177717
rect 107028 177712 107627 177714
rect 107028 177656 107566 177712
rect 107622 177656 107627 177712
rect 107028 177654 107627 177656
rect 107028 177652 107034 177654
rect 107561 177651 107627 177654
rect 114318 177652 114324 177716
rect 114388 177714 114394 177716
rect 114461 177714 114527 177717
rect 116945 177716 117011 177717
rect 116894 177714 116900 177716
rect 114388 177712 114527 177714
rect 114388 177656 114466 177712
rect 114522 177656 114527 177712
rect 114388 177654 114527 177656
rect 116854 177654 116900 177714
rect 116964 177712 117011 177716
rect 117006 177656 117011 177712
rect 114388 177652 114394 177654
rect 114461 177651 114527 177654
rect 116894 177652 116900 177654
rect 116964 177652 117011 177656
rect 118366 177652 118372 177716
rect 118436 177714 118442 177716
rect 118601 177714 118667 177717
rect 118436 177712 118667 177714
rect 118436 177656 118606 177712
rect 118662 177656 118667 177712
rect 118436 177654 118667 177656
rect 118436 177652 118442 177654
rect 116945 177651 117011 177652
rect 118601 177651 118667 177654
rect 120758 177652 120764 177716
rect 120828 177714 120834 177716
rect 121361 177714 121427 177717
rect 129457 177716 129523 177717
rect 132401 177716 132467 177717
rect 129406 177714 129412 177716
rect 120828 177712 121427 177714
rect 120828 177656 121366 177712
rect 121422 177656 121427 177712
rect 120828 177654 121427 177656
rect 129366 177654 129412 177714
rect 129476 177712 129523 177716
rect 132350 177714 132356 177716
rect 129518 177656 129523 177712
rect 120828 177652 120834 177654
rect 121361 177651 121427 177654
rect 129406 177652 129412 177654
rect 129476 177652 129523 177656
rect 132310 177654 132356 177714
rect 132420 177712 132467 177716
rect 132462 177656 132467 177712
rect 132350 177652 132356 177654
rect 132420 177652 132467 177656
rect 133086 177652 133092 177716
rect 133156 177714 133162 177716
rect 133781 177714 133847 177717
rect 133156 177712 133847 177714
rect 133156 177656 133786 177712
rect 133842 177656 133847 177712
rect 133156 177654 133847 177656
rect 133156 177652 133162 177654
rect 129457 177651 129523 177652
rect 132401 177651 132467 177652
rect 133781 177651 133847 177654
rect 232497 177578 232563 177581
rect 258390 177578 258396 177580
rect 232497 177576 258396 177578
rect 232497 177520 232502 177576
rect 232558 177520 258396 177576
rect 232497 177518 258396 177520
rect 232497 177515 232563 177518
rect 258390 177516 258396 177518
rect 258460 177516 258466 177580
rect 226977 177442 227043 177445
rect 259494 177442 259500 177444
rect 226977 177440 259500 177442
rect 226977 177384 226982 177440
rect 227038 177384 259500 177440
rect 226977 177382 259500 177384
rect 226977 177379 227043 177382
rect 259494 177380 259500 177382
rect 259564 177380 259570 177444
rect 178677 177306 178743 177309
rect 249374 177306 249380 177308
rect 178677 177304 249380 177306
rect 178677 177248 178682 177304
rect 178738 177248 249380 177304
rect 178677 177246 249380 177248
rect 178677 177243 178743 177246
rect 249374 177244 249380 177246
rect 249444 177244 249450 177308
rect 286317 177306 286383 177309
rect 331438 177306 331444 177308
rect 286317 177304 331444 177306
rect 286317 177248 286322 177304
rect 286378 177248 331444 177304
rect 286317 177246 331444 177248
rect 286317 177243 286383 177246
rect 331438 177244 331444 177246
rect 331508 177244 331514 177308
rect 112110 177108 112116 177172
rect 112180 177170 112186 177172
rect 112989 177170 113055 177173
rect 112180 177168 113055 177170
rect 112180 177112 112994 177168
rect 113050 177112 113055 177168
rect 112180 177110 113055 177112
rect 112180 177108 112186 177110
rect 112989 177107 113055 177110
rect 110689 177036 110755 177037
rect 110638 177034 110644 177036
rect 110598 176974 110644 177034
rect 110708 177032 110755 177036
rect 110750 176976 110755 177032
rect 110638 176972 110644 176974
rect 110708 176972 110755 176976
rect 123150 176972 123156 177036
rect 123220 177034 123226 177036
rect 123753 177034 123819 177037
rect 123220 177032 123819 177034
rect 123220 176976 123758 177032
rect 123814 176976 123819 177032
rect 123220 176974 123819 176976
rect 123220 176972 123226 176974
rect 110689 176971 110755 176972
rect 123753 176971 123819 176974
rect 127014 176972 127020 177036
rect 127084 177034 127090 177036
rect 128077 177034 128143 177037
rect 127084 177032 128143 177034
rect 127084 176976 128082 177032
rect 128138 176976 128143 177032
rect 127084 176974 128143 176976
rect 127084 176972 127090 176974
rect 128077 176971 128143 176974
rect 101990 176836 101996 176900
rect 102060 176898 102066 176900
rect 186957 176898 187023 176901
rect 102060 176896 187023 176898
rect 102060 176840 186962 176896
rect 187018 176840 187023 176896
rect 102060 176838 187023 176840
rect 102060 176836 102066 176838
rect 186957 176835 187023 176838
rect 100661 176762 100727 176765
rect 103329 176762 103395 176765
rect 104617 176764 104683 176765
rect 108113 176764 108179 176765
rect 104566 176762 104572 176764
rect 99422 176760 100727 176762
rect 99422 176704 100666 176760
rect 100722 176704 100727 176760
rect 99422 176702 100727 176704
rect 99422 176492 99482 176702
rect 100661 176699 100727 176702
rect 103286 176760 103395 176762
rect 103286 176704 103334 176760
rect 103390 176704 103395 176760
rect 103286 176699 103395 176704
rect 104526 176702 104572 176762
rect 104636 176760 104683 176764
rect 108062 176762 108068 176764
rect 104678 176704 104683 176760
rect 104566 176700 104572 176702
rect 104636 176700 104683 176704
rect 108022 176702 108068 176762
rect 108132 176760 108179 176764
rect 108174 176704 108179 176760
rect 108062 176700 108068 176702
rect 108132 176700 108179 176704
rect 109534 176700 109540 176764
rect 109604 176762 109610 176764
rect 109953 176762 110019 176765
rect 115841 176764 115907 176765
rect 124489 176764 124555 176765
rect 115790 176762 115796 176764
rect 109604 176760 110019 176762
rect 109604 176704 109958 176760
rect 110014 176704 110019 176760
rect 109604 176702 110019 176704
rect 115750 176702 115796 176762
rect 115860 176760 115907 176764
rect 124438 176762 124444 176764
rect 115902 176704 115907 176760
rect 109604 176700 109610 176702
rect 104617 176699 104683 176700
rect 108113 176699 108179 176700
rect 109953 176699 110019 176702
rect 115790 176700 115796 176702
rect 115860 176700 115907 176704
rect 124398 176702 124444 176762
rect 124508 176760 124555 176764
rect 124550 176704 124555 176760
rect 124438 176700 124444 176702
rect 124508 176700 124555 176704
rect 125726 176700 125732 176764
rect 125796 176762 125802 176764
rect 126053 176762 126119 176765
rect 130745 176764 130811 176765
rect 130694 176762 130700 176764
rect 125796 176760 126119 176762
rect 125796 176704 126058 176760
rect 126114 176704 126119 176760
rect 125796 176702 126119 176704
rect 130654 176702 130700 176762
rect 130764 176760 130811 176764
rect 130806 176704 130811 176760
rect 125796 176700 125802 176702
rect 115841 176699 115907 176700
rect 124489 176699 124555 176700
rect 126053 176699 126119 176702
rect 130694 176700 130700 176702
rect 130764 176700 130811 176704
rect 134374 176700 134380 176764
rect 134444 176762 134450 176764
rect 134793 176762 134859 176765
rect 136081 176764 136147 176765
rect 148225 176764 148291 176765
rect 136030 176762 136036 176764
rect 134444 176760 134859 176762
rect 134444 176704 134798 176760
rect 134854 176704 134859 176760
rect 134444 176702 134859 176704
rect 135990 176702 136036 176762
rect 136100 176760 136147 176764
rect 148174 176762 148180 176764
rect 136142 176704 136147 176760
rect 134444 176700 134450 176702
rect 130745 176699 130811 176700
rect 134793 176699 134859 176702
rect 136030 176700 136036 176702
rect 136100 176700 136147 176704
rect 148134 176702 148180 176762
rect 148244 176760 148291 176764
rect 148286 176704 148291 176760
rect 148174 176700 148180 176702
rect 148244 176700 148291 176704
rect 260046 176700 260052 176764
rect 260116 176762 260122 176764
rect 316033 176762 316099 176765
rect 260116 176760 316099 176762
rect 260116 176704 316038 176760
rect 316094 176704 316099 176760
rect 260116 176702 316099 176704
rect 260116 176700 260122 176702
rect 136081 176699 136147 176700
rect 148225 176699 148291 176700
rect 316033 176699 316099 176702
rect 103286 176492 103346 176699
rect 99414 176428 99420 176492
rect 99484 176428 99490 176492
rect 103278 176428 103284 176492
rect 103348 176428 103354 176492
rect 213913 176218 213979 176221
rect 316309 176218 316375 176221
rect 213913 176216 217242 176218
rect 213913 176160 213918 176216
rect 213974 176160 217242 176216
rect 213913 176158 217242 176160
rect 213913 176155 213979 176158
rect -960 175796 480 176036
rect 217182 175644 217242 176158
rect 316309 176216 325710 176218
rect 316309 176160 316314 176216
rect 316370 176160 325710 176216
rect 316309 176158 325710 176160
rect 316309 176155 316375 176158
rect 224217 176082 224283 176085
rect 249190 176082 249196 176084
rect 224217 176080 249196 176082
rect 224217 176024 224222 176080
rect 224278 176024 249196 176080
rect 224217 176022 249196 176024
rect 224217 176019 224283 176022
rect 249190 176020 249196 176022
rect 249260 176020 249266 176084
rect 321461 176082 321527 176085
rect 321461 176080 321570 176082
rect 321461 176024 321466 176080
rect 321522 176024 321570 176080
rect 321461 176019 321570 176024
rect 220077 175946 220143 175949
rect 260966 175946 260972 175948
rect 220077 175944 260972 175946
rect 220077 175888 220082 175944
rect 220138 175888 260972 175944
rect 220077 175886 260972 175888
rect 220077 175883 220143 175886
rect 260966 175884 260972 175886
rect 261036 175884 261042 175948
rect 246941 175810 247007 175813
rect 246941 175808 248338 175810
rect 246941 175752 246946 175808
rect 247002 175752 248338 175808
rect 246941 175750 248338 175752
rect 246941 175747 247007 175750
rect 248278 175644 248338 175750
rect 296670 175614 310132 175674
rect 100753 175404 100819 175405
rect 121913 175404 121979 175405
rect 128169 175404 128235 175405
rect 158897 175404 158963 175405
rect 100702 175402 100708 175404
rect 100662 175342 100708 175402
rect 100772 175400 100819 175404
rect 121862 175402 121868 175404
rect 100814 175344 100819 175400
rect 100702 175340 100708 175342
rect 100772 175340 100819 175344
rect 121822 175342 121868 175402
rect 121932 175400 121979 175404
rect 128118 175402 128124 175404
rect 121974 175344 121979 175400
rect 121862 175340 121868 175342
rect 121932 175340 121979 175344
rect 128078 175342 128124 175402
rect 128188 175400 128235 175404
rect 158846 175402 158852 175404
rect 128230 175344 128235 175400
rect 128118 175340 128124 175342
rect 128188 175340 128235 175344
rect 158806 175342 158852 175402
rect 158916 175400 158963 175404
rect 158958 175344 158963 175400
rect 158846 175340 158852 175342
rect 158916 175340 158963 175344
rect 262806 175340 262812 175404
rect 262876 175402 262882 175404
rect 296670 175402 296730 175614
rect 321510 175508 321570 176019
rect 325650 175946 325710 176158
rect 325969 175946 326035 175949
rect 325650 175944 326035 175946
rect 325650 175888 325974 175944
rect 326030 175888 326035 175944
rect 325650 175886 326035 175888
rect 325969 175883 326035 175886
rect 262876 175342 296730 175402
rect 262876 175340 262882 175342
rect 100753 175339 100819 175340
rect 121913 175339 121979 175340
rect 128169 175339 128235 175340
rect 158897 175339 158963 175340
rect 249241 175266 249307 175269
rect 248952 175264 249307 175266
rect 248952 175208 249246 175264
rect 249302 175208 249307 175264
rect 248952 175206 249307 175208
rect 249241 175203 249307 175206
rect 307109 175266 307175 175269
rect 321461 175266 321527 175269
rect 307109 175264 310040 175266
rect 307109 175208 307114 175264
rect 307170 175208 310040 175264
rect 307109 175206 310040 175208
rect 321461 175264 321570 175266
rect 321461 175208 321466 175264
rect 321522 175208 321570 175264
rect 307109 175203 307175 175206
rect 321461 175203 321570 175208
rect 213913 175130 213979 175133
rect 213913 175128 217242 175130
rect 213913 175072 213918 175128
rect 213974 175072 217242 175128
rect 213913 175070 217242 175072
rect 213913 175067 213979 175070
rect 113173 174996 113239 174997
rect 119429 174996 119495 174997
rect 113136 174932 113142 174996
rect 113206 174994 113239 174996
rect 119392 174994 119398 174996
rect 113206 174992 113298 174994
rect 113234 174936 113298 174992
rect 113206 174934 113298 174936
rect 119338 174934 119398 174994
rect 119462 174992 119495 174996
rect 119490 174936 119495 174992
rect 217182 174964 217242 175070
rect 113206 174932 113239 174934
rect 119392 174932 119398 174934
rect 119462 174932 119495 174936
rect 113173 174931 113239 174932
rect 119429 174931 119495 174932
rect 306557 174858 306623 174861
rect 306557 174856 310040 174858
rect 306557 174800 306562 174856
rect 306618 174800 310040 174856
rect 306557 174798 310040 174800
rect 306557 174795 306623 174798
rect 214557 174722 214623 174725
rect 249149 174722 249215 174725
rect 214557 174720 217242 174722
rect 214557 174664 214562 174720
rect 214618 174664 217242 174720
rect 214557 174662 217242 174664
rect 248952 174720 249215 174722
rect 248952 174664 249154 174720
rect 249210 174664 249215 174720
rect 321510 174692 321570 175203
rect 248952 174662 249215 174664
rect 214557 174659 214623 174662
rect 217182 174284 217242 174662
rect 249149 174659 249215 174662
rect 307569 174450 307635 174453
rect 307569 174448 310040 174450
rect 307569 174392 307574 174448
rect 307630 174392 310040 174448
rect 307569 174390 310040 174392
rect 307569 174387 307635 174390
rect 249190 174314 249196 174316
rect 248952 174254 249196 174314
rect 249190 174252 249196 174254
rect 249260 174252 249266 174316
rect 307661 174042 307727 174045
rect 324497 174042 324563 174045
rect 307661 174040 310040 174042
rect 307661 173984 307666 174040
rect 307722 173984 310040 174040
rect 307661 173982 310040 173984
rect 321908 174040 324563 174042
rect 321908 173984 324502 174040
rect 324558 173984 324563 174040
rect 321908 173982 324563 173984
rect 307661 173979 307727 173982
rect 324497 173979 324563 173982
rect 213913 173770 213979 173773
rect 252461 173770 252527 173773
rect 213913 173768 217242 173770
rect 213913 173712 213918 173768
rect 213974 173712 217242 173768
rect 213913 173710 217242 173712
rect 248952 173768 252527 173770
rect 248952 173712 252466 173768
rect 252522 173712 252527 173768
rect 248952 173710 252527 173712
rect 213913 173707 213979 173710
rect 217182 173604 217242 173710
rect 252461 173707 252527 173710
rect 307569 173634 307635 173637
rect 307569 173632 310040 173634
rect 307569 173576 307574 173632
rect 307630 173576 310040 173632
rect 307569 173574 310040 173576
rect 307569 173571 307635 173574
rect 214005 173362 214071 173365
rect 249374 173362 249380 173364
rect 214005 173360 217242 173362
rect 214005 173304 214010 173360
rect 214066 173304 217242 173360
rect 214005 173302 217242 173304
rect 248952 173302 249380 173362
rect 214005 173299 214071 173302
rect 217182 172924 217242 173302
rect 249374 173300 249380 173302
rect 249444 173300 249450 173364
rect 307661 173226 307727 173229
rect 324589 173226 324655 173229
rect 307661 173224 310040 173226
rect 307661 173168 307666 173224
rect 307722 173168 310040 173224
rect 307661 173166 310040 173168
rect 321908 173224 324655 173226
rect 321908 173168 324594 173224
rect 324650 173168 324655 173224
rect 321908 173166 324655 173168
rect 307661 173163 307727 173166
rect 324589 173163 324655 173166
rect 249149 172802 249215 172805
rect 248860 172800 249215 172802
rect 248860 172744 249154 172800
rect 249210 172744 249215 172800
rect 248860 172742 249215 172744
rect 249149 172739 249215 172742
rect 307477 172682 307543 172685
rect 307477 172680 310040 172682
rect 307477 172624 307482 172680
rect 307538 172624 310040 172680
rect 307477 172622 310040 172624
rect 307477 172619 307543 172622
rect 213269 172410 213335 172413
rect 252369 172410 252435 172413
rect 324313 172410 324379 172413
rect 213269 172408 217242 172410
rect 213269 172352 213274 172408
rect 213330 172352 217242 172408
rect 213269 172350 217242 172352
rect 248952 172408 252435 172410
rect 248952 172352 252374 172408
rect 252430 172352 252435 172408
rect 248952 172350 252435 172352
rect 321908 172408 324379 172410
rect 321908 172352 324318 172408
rect 324374 172352 324379 172408
rect 321908 172350 324379 172352
rect 213269 172347 213335 172350
rect 217182 172244 217242 172350
rect 252369 172347 252435 172350
rect 324313 172347 324379 172350
rect 306557 172274 306623 172277
rect 306557 172272 310040 172274
rect 306557 172216 306562 172272
rect 306618 172216 310040 172272
rect 306557 172214 310040 172216
rect 306557 172211 306623 172214
rect 213913 172002 213979 172005
rect 213913 172000 217242 172002
rect 213913 171944 213918 172000
rect 213974 171944 217242 172000
rect 213913 171942 217242 171944
rect 213913 171939 213979 171942
rect 168005 171594 168071 171597
rect 164694 171592 168071 171594
rect 164694 171536 168010 171592
rect 168066 171536 168071 171592
rect 217182 171564 217242 171942
rect 252645 171866 252711 171869
rect 248952 171864 252711 171866
rect 248952 171808 252650 171864
rect 252706 171808 252711 171864
rect 248952 171806 252711 171808
rect 252645 171803 252711 171806
rect 307569 171866 307635 171869
rect 307569 171864 310040 171866
rect 307569 171808 307574 171864
rect 307630 171808 310040 171864
rect 307569 171806 310040 171808
rect 307569 171803 307635 171806
rect 164694 171534 168071 171536
rect 168005 171531 168071 171534
rect 252461 171458 252527 171461
rect 248952 171456 252527 171458
rect 248952 171400 252466 171456
rect 252522 171400 252527 171456
rect 248952 171398 252527 171400
rect 252461 171395 252527 171398
rect 307661 171458 307727 171461
rect 307661 171456 310040 171458
rect 307661 171400 307666 171456
rect 307722 171400 310040 171456
rect 307661 171398 310040 171400
rect 307661 171395 307727 171398
rect 321878 171186 321938 171700
rect 325969 171186 326035 171189
rect 216998 171126 217242 171186
rect 321878 171184 326035 171186
rect 321878 171128 325974 171184
rect 326030 171128 326035 171184
rect 321878 171126 326035 171128
rect 216998 171050 217058 171126
rect 215250 170990 217058 171050
rect 217182 171020 217242 171126
rect 325969 171123 326035 171126
rect 307569 171050 307635 171053
rect 307569 171048 310040 171050
rect 307569 170992 307574 171048
rect 307630 170992 310040 171048
rect 307569 170990 310040 170992
rect 214465 170914 214531 170917
rect 215250 170914 215310 170990
rect 307569 170987 307635 170990
rect 324313 170914 324379 170917
rect 214465 170912 215310 170914
rect 214465 170856 214470 170912
rect 214526 170856 215310 170912
rect 321908 170912 324379 170914
rect 214465 170854 215310 170856
rect 214465 170851 214531 170854
rect 248860 170810 249442 170870
rect 321908 170856 324318 170912
rect 324374 170856 324379 170912
rect 321908 170854 324379 170856
rect 324313 170851 324379 170854
rect 213913 170778 213979 170781
rect 213913 170776 217242 170778
rect 213913 170720 213918 170776
rect 213974 170720 217242 170776
rect 213913 170718 217242 170720
rect 213913 170715 213979 170718
rect 217182 170340 217242 170718
rect 248860 170402 249258 170462
rect 249198 170234 249258 170402
rect 249382 170370 249442 170810
rect 306557 170642 306623 170645
rect 306557 170640 310040 170642
rect 306557 170584 306562 170640
rect 306618 170584 310040 170640
rect 306557 170582 310040 170584
rect 306557 170579 306623 170582
rect 321318 170580 321324 170644
rect 321388 170580 321394 170644
rect 260966 170370 260972 170372
rect 249382 170310 260972 170370
rect 260966 170308 260972 170310
rect 261036 170308 261042 170372
rect 252461 170234 252527 170237
rect 249198 170232 252527 170234
rect 249198 170176 252466 170232
rect 252522 170176 252527 170232
rect 249198 170174 252527 170176
rect 252461 170171 252527 170174
rect 307661 170234 307727 170237
rect 307661 170232 310040 170234
rect 307661 170176 307666 170232
rect 307722 170176 310040 170232
rect 307661 170174 310040 170176
rect 307661 170171 307727 170174
rect 252461 170098 252527 170101
rect 248952 170096 252527 170098
rect 248952 170040 252466 170096
rect 252522 170040 252527 170096
rect 321326 170068 321386 170580
rect 248952 170038 252527 170040
rect 252461 170035 252527 170038
rect 307385 169826 307451 169829
rect 216998 169766 217242 169826
rect 214005 169690 214071 169693
rect 216998 169690 217058 169766
rect 214005 169688 217058 169690
rect 214005 169632 214010 169688
rect 214066 169632 217058 169688
rect 217182 169660 217242 169766
rect 307385 169824 310040 169826
rect 307385 169768 307390 169824
rect 307446 169768 310040 169824
rect 307385 169766 310040 169768
rect 307385 169763 307451 169766
rect 321277 169690 321343 169693
rect 321277 169688 321386 169690
rect 214005 169630 217058 169632
rect 321277 169632 321282 169688
rect 321338 169632 321386 169688
rect 214005 169627 214071 169630
rect 321277 169627 321386 169632
rect 252461 169554 252527 169557
rect 248952 169552 252527 169554
rect 248952 169496 252466 169552
rect 252522 169496 252527 169552
rect 248952 169494 252527 169496
rect 252461 169491 252527 169494
rect 213913 169418 213979 169421
rect 213913 169416 217242 169418
rect 213913 169360 213918 169416
rect 213974 169360 217242 169416
rect 321326 169388 321386 169627
rect 213913 169358 217242 169360
rect 213913 169355 213979 169358
rect 217182 168980 217242 169358
rect 307661 169282 307727 169285
rect 307661 169280 310040 169282
rect 307661 169224 307666 169280
rect 307722 169224 310040 169280
rect 307661 169222 310040 169224
rect 307661 169219 307727 169222
rect 252369 169146 252435 169149
rect 248952 169144 252435 169146
rect 248952 169088 252374 169144
rect 252430 169088 252435 169144
rect 248952 169086 252435 169088
rect 252369 169083 252435 169086
rect 307569 168874 307635 168877
rect 307569 168872 310040 168874
rect 307569 168816 307574 168872
rect 307630 168816 310040 168872
rect 307569 168814 310040 168816
rect 307569 168811 307635 168814
rect 252277 168602 252343 168605
rect 324405 168602 324471 168605
rect 248952 168600 252343 168602
rect 248952 168544 252282 168600
rect 252338 168544 252343 168600
rect 248952 168542 252343 168544
rect 321908 168600 324471 168602
rect 321908 168544 324410 168600
rect 324466 168544 324471 168600
rect 321908 168542 324471 168544
rect 252277 168539 252343 168542
rect 324405 168539 324471 168542
rect 307477 168466 307543 168469
rect 307477 168464 310040 168466
rect 307477 168408 307482 168464
rect 307538 168408 310040 168464
rect 307477 168406 310040 168408
rect 307477 168403 307543 168406
rect 213913 168058 213979 168061
rect 217182 168058 217242 168300
rect 252461 168194 252527 168197
rect 248952 168192 252527 168194
rect 248952 168136 252466 168192
rect 252522 168136 252527 168192
rect 248952 168134 252527 168136
rect 252461 168131 252527 168134
rect 213913 168056 217242 168058
rect 213913 168000 213918 168056
rect 213974 168000 217242 168056
rect 213913 167998 217242 168000
rect 307477 168058 307543 168061
rect 307477 168056 310040 168058
rect 307477 168000 307482 168056
rect 307538 168000 310040 168056
rect 307477 167998 310040 168000
rect 213913 167995 213979 167998
rect 307477 167995 307543 167998
rect 214005 167922 214071 167925
rect 214005 167920 217242 167922
rect 214005 167864 214010 167920
rect 214066 167864 217242 167920
rect 214005 167862 217242 167864
rect 214005 167859 214071 167862
rect 217182 167620 217242 167862
rect 324313 167786 324379 167789
rect 321908 167784 324379 167786
rect 321908 167728 324318 167784
rect 324374 167728 324379 167784
rect 321908 167726 324379 167728
rect 324313 167723 324379 167726
rect 252277 167650 252343 167653
rect 248952 167648 252343 167650
rect 248952 167592 252282 167648
rect 252338 167592 252343 167648
rect 248952 167590 252343 167592
rect 252277 167587 252343 167590
rect 307569 167650 307635 167653
rect 307569 167648 310040 167650
rect 307569 167592 307574 167648
rect 307630 167592 310040 167648
rect 307569 167590 310040 167592
rect 307569 167587 307635 167590
rect 252369 167242 252435 167245
rect 248952 167240 252435 167242
rect 248952 167184 252374 167240
rect 252430 167184 252435 167240
rect 248952 167182 252435 167184
rect 252369 167179 252435 167182
rect 307661 167242 307727 167245
rect 307661 167240 310040 167242
rect 307661 167184 307666 167240
rect 307722 167184 310040 167240
rect 307661 167182 310040 167184
rect 307661 167179 307727 167182
rect 324405 167106 324471 167109
rect 321908 167104 324471 167106
rect 321908 167048 324410 167104
rect 324466 167048 324471 167104
rect 321908 167046 324471 167048
rect 324405 167043 324471 167046
rect 214741 166970 214807 166973
rect 216998 166970 217242 167010
rect 214741 166968 217242 166970
rect 214741 166912 214746 166968
rect 214802 166950 217242 166968
rect 214802 166912 217058 166950
rect 217182 166940 217242 166950
rect 214741 166910 217058 166912
rect 214741 166907 214807 166910
rect 307569 166834 307635 166837
rect 307569 166832 310040 166834
rect 307569 166776 307574 166832
rect 307630 166776 310040 166832
rect 307569 166774 310040 166776
rect 307569 166771 307635 166774
rect 214465 166698 214531 166701
rect 252461 166698 252527 166701
rect 214465 166696 217242 166698
rect 214465 166640 214470 166696
rect 214526 166640 217242 166696
rect 214465 166638 217242 166640
rect 248952 166696 252527 166698
rect 248952 166640 252466 166696
rect 252522 166640 252527 166696
rect 248952 166638 252527 166640
rect 214465 166635 214531 166638
rect 217182 166396 217242 166638
rect 252461 166635 252527 166638
rect 307293 166426 307359 166429
rect 307293 166424 310040 166426
rect 307293 166368 307298 166424
rect 307354 166368 310040 166424
rect 307293 166366 310040 166368
rect 307293 166363 307359 166366
rect 252369 166290 252435 166293
rect 324313 166290 324379 166293
rect 248952 166288 252435 166290
rect 248952 166232 252374 166288
rect 252430 166232 252435 166288
rect 248952 166230 252435 166232
rect 321908 166288 324379 166290
rect 321908 166232 324318 166288
rect 324374 166232 324379 166288
rect 321908 166230 324379 166232
rect 252369 166227 252435 166230
rect 324313 166227 324379 166230
rect 213913 166154 213979 166157
rect 213913 166152 217242 166154
rect 213913 166096 213918 166152
rect 213974 166096 217242 166152
rect 213913 166094 217242 166096
rect 213913 166091 213979 166094
rect 217182 165716 217242 166094
rect 307661 165882 307727 165885
rect 583520 165882 584960 165972
rect 307661 165880 310040 165882
rect 307661 165824 307666 165880
rect 307722 165824 310040 165880
rect 307661 165822 310040 165824
rect 567150 165822 584960 165882
rect 307661 165819 307727 165822
rect 249885 165746 249951 165749
rect 248952 165744 249951 165746
rect 248952 165688 249890 165744
rect 249946 165688 249951 165744
rect 248952 165686 249951 165688
rect 249885 165683 249951 165686
rect 338614 165684 338620 165748
rect 338684 165746 338690 165748
rect 567150 165746 567210 165822
rect 338684 165686 567210 165746
rect 583520 165732 584960 165822
rect 338684 165684 338690 165686
rect 307293 165474 307359 165477
rect 323209 165474 323275 165477
rect 307293 165472 310040 165474
rect 307293 165416 307298 165472
rect 307354 165416 310040 165472
rect 307293 165414 310040 165416
rect 321908 165472 323275 165474
rect 321908 165416 323214 165472
rect 323270 165416 323275 165472
rect 321908 165414 323275 165416
rect 307293 165411 307359 165414
rect 323209 165411 323275 165414
rect 213913 165338 213979 165341
rect 252461 165338 252527 165341
rect 213913 165336 217242 165338
rect 213913 165280 213918 165336
rect 213974 165280 217242 165336
rect 213913 165278 217242 165280
rect 248952 165336 252527 165338
rect 248952 165280 252466 165336
rect 252522 165280 252527 165336
rect 248952 165278 252527 165280
rect 213913 165275 213979 165278
rect 217182 165036 217242 165278
rect 252461 165275 252527 165278
rect 307017 165066 307083 165069
rect 307017 165064 310040 165066
rect 307017 165008 307022 165064
rect 307078 165008 310040 165064
rect 307017 165006 310040 165008
rect 307017 165003 307083 165006
rect 214005 164794 214071 164797
rect 252369 164794 252435 164797
rect 324313 164794 324379 164797
rect 214005 164792 217242 164794
rect 214005 164736 214010 164792
rect 214066 164736 217242 164792
rect 214005 164734 217242 164736
rect 248952 164792 252435 164794
rect 248952 164736 252374 164792
rect 252430 164736 252435 164792
rect 248952 164734 252435 164736
rect 321908 164792 324379 164794
rect 321908 164736 324318 164792
rect 324374 164736 324379 164792
rect 321908 164734 324379 164736
rect 214005 164731 214071 164734
rect 217182 164356 217242 164734
rect 252369 164731 252435 164734
rect 324313 164731 324379 164734
rect 307661 164658 307727 164661
rect 307661 164656 310040 164658
rect 307661 164600 307666 164656
rect 307722 164600 310040 164656
rect 307661 164598 310040 164600
rect 307661 164595 307727 164598
rect 252737 164386 252803 164389
rect 248952 164384 252803 164386
rect 248952 164328 252742 164384
rect 252798 164328 252803 164384
rect 248952 164326 252803 164328
rect 252737 164323 252803 164326
rect 307569 164250 307635 164253
rect 307569 164248 310040 164250
rect 307569 164192 307574 164248
rect 307630 164192 310040 164248
rect 307569 164190 310040 164192
rect 307569 164187 307635 164190
rect 213913 164114 213979 164117
rect 213913 164112 217242 164114
rect 213913 164056 213918 164112
rect 213974 164056 217242 164112
rect 213913 164054 217242 164056
rect 213913 164051 213979 164054
rect 217182 163676 217242 164054
rect 252461 163978 252527 163981
rect 324313 163978 324379 163981
rect 248952 163976 252527 163978
rect 248952 163920 252466 163976
rect 252522 163920 252527 163976
rect 248952 163918 252527 163920
rect 321908 163976 324379 163978
rect 321908 163920 324318 163976
rect 324374 163920 324379 163976
rect 321908 163918 324379 163920
rect 252461 163915 252527 163918
rect 324313 163915 324379 163918
rect 307569 163842 307635 163845
rect 307569 163840 310040 163842
rect 307569 163784 307574 163840
rect 307630 163784 310040 163840
rect 307569 163782 310040 163784
rect 307569 163779 307635 163782
rect 214005 163434 214071 163437
rect 254526 163434 254532 163436
rect 214005 163432 217242 163434
rect 214005 163376 214010 163432
rect 214066 163376 217242 163432
rect 214005 163374 217242 163376
rect 248952 163374 254532 163434
rect 214005 163371 214071 163374
rect 217182 162996 217242 163374
rect 254526 163372 254532 163374
rect 254596 163372 254602 163436
rect 307477 163434 307543 163437
rect 307477 163432 310040 163434
rect 307477 163376 307482 163432
rect 307538 163376 310040 163432
rect 307477 163374 310040 163376
rect 307477 163371 307543 163374
rect 324405 163162 324471 163165
rect 321908 163160 324471 163162
rect 321908 163104 324410 163160
rect 324466 163104 324471 163160
rect 321908 163102 324471 163104
rect 324405 163099 324471 163102
rect 251449 163026 251515 163029
rect 248952 163024 251515 163026
rect -960 162890 480 162980
rect 248952 162968 251454 163024
rect 251510 162968 251515 163024
rect 248952 162966 251515 162968
rect 251449 162963 251515 162966
rect 307661 163026 307727 163029
rect 307661 163024 310040 163026
rect 307661 162968 307666 163024
rect 307722 162968 310040 163024
rect 307661 162966 310040 162968
rect 307661 162963 307727 162966
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 252461 162482 252527 162485
rect 248952 162480 252527 162482
rect 248952 162424 252466 162480
rect 252522 162424 252527 162480
rect 248952 162422 252527 162424
rect 252461 162419 252527 162422
rect 307569 162482 307635 162485
rect 324313 162482 324379 162485
rect 307569 162480 310040 162482
rect 307569 162424 307574 162480
rect 307630 162424 310040 162480
rect 307569 162422 310040 162424
rect 321908 162480 324379 162482
rect 321908 162424 324318 162480
rect 324374 162424 324379 162480
rect 321908 162422 324379 162424
rect 307569 162419 307635 162422
rect 324313 162419 324379 162422
rect 217182 161938 217242 162316
rect 252369 162074 252435 162077
rect 248952 162072 252435 162074
rect 248952 162016 252374 162072
rect 252430 162016 252435 162072
rect 248952 162014 252435 162016
rect 252369 162011 252435 162014
rect 307477 162074 307543 162077
rect 307477 162072 310040 162074
rect 307477 162016 307482 162072
rect 307538 162016 310040 162072
rect 307477 162014 310040 162016
rect 307477 162011 307543 162014
rect 200070 161878 217242 161938
rect 166390 161468 166396 161532
rect 166460 161530 166466 161532
rect 200070 161530 200130 161878
rect 166460 161470 200130 161530
rect 213913 161530 213979 161533
rect 217366 161530 217426 161772
rect 307661 161666 307727 161669
rect 324313 161666 324379 161669
rect 307661 161664 310040 161666
rect 307661 161608 307666 161664
rect 307722 161608 310040 161664
rect 307661 161606 310040 161608
rect 321908 161664 324379 161666
rect 321908 161608 324318 161664
rect 324374 161608 324379 161664
rect 321908 161606 324379 161608
rect 307661 161603 307727 161606
rect 324313 161603 324379 161606
rect 252277 161530 252343 161533
rect 213913 161528 217426 161530
rect 213913 161472 213918 161528
rect 213974 161472 217426 161528
rect 213913 161470 217426 161472
rect 248952 161528 252343 161530
rect 248952 161472 252282 161528
rect 252338 161472 252343 161528
rect 248952 161470 252343 161472
rect 166460 161468 166466 161470
rect 213913 161467 213979 161470
rect 252277 161467 252343 161470
rect 213913 161258 213979 161261
rect 307569 161258 307635 161261
rect 213913 161256 217242 161258
rect 213913 161200 213918 161256
rect 213974 161200 217242 161256
rect 213913 161198 217242 161200
rect 213913 161195 213979 161198
rect 217182 161092 217242 161198
rect 307569 161256 310040 161258
rect 307569 161200 307574 161256
rect 307630 161200 310040 161256
rect 307569 161198 310040 161200
rect 307569 161195 307635 161198
rect 248860 161018 249442 161078
rect 214005 160850 214071 160853
rect 249382 160850 249442 161018
rect 259494 160850 259500 160852
rect 214005 160848 217242 160850
rect 214005 160792 214010 160848
rect 214066 160792 217242 160848
rect 214005 160790 217242 160792
rect 249382 160790 259500 160850
rect 214005 160787 214071 160790
rect 217182 160412 217242 160790
rect 259494 160788 259500 160790
rect 259564 160788 259570 160852
rect 307201 160850 307267 160853
rect 324313 160850 324379 160853
rect 307201 160848 310040 160850
rect 307201 160792 307206 160848
rect 307262 160792 310040 160848
rect 307201 160790 310040 160792
rect 321908 160848 324379 160850
rect 321908 160792 324318 160848
rect 324374 160792 324379 160848
rect 321908 160790 324379 160792
rect 307201 160787 307267 160790
rect 324313 160787 324379 160790
rect 252461 160578 252527 160581
rect 248952 160576 252527 160578
rect 248952 160520 252466 160576
rect 252522 160520 252527 160576
rect 248952 160518 252527 160520
rect 252461 160515 252527 160518
rect 307661 160442 307727 160445
rect 307661 160440 310040 160442
rect 307661 160384 307666 160440
rect 307722 160384 310040 160440
rect 307661 160382 310040 160384
rect 307661 160379 307727 160382
rect 251357 160170 251423 160173
rect 324405 160170 324471 160173
rect 248952 160168 251423 160170
rect 248952 160112 251362 160168
rect 251418 160112 251423 160168
rect 248952 160110 251423 160112
rect 321908 160168 324471 160170
rect 321908 160112 324410 160168
rect 324466 160112 324471 160168
rect 321908 160110 324471 160112
rect 251357 160107 251423 160110
rect 324405 160107 324471 160110
rect 213913 160034 213979 160037
rect 307293 160034 307359 160037
rect 213913 160032 217242 160034
rect 213913 159976 213918 160032
rect 213974 159976 217242 160032
rect 213913 159974 217242 159976
rect 213913 159971 213979 159974
rect 217182 159732 217242 159974
rect 307293 160032 310040 160034
rect 307293 159976 307298 160032
rect 307354 159976 310040 160032
rect 307293 159974 310040 159976
rect 307293 159971 307359 159974
rect 252461 159626 252527 159629
rect 248952 159624 252527 159626
rect 248952 159568 252466 159624
rect 252522 159568 252527 159624
rect 248952 159566 252527 159568
rect 252461 159563 252527 159566
rect 307661 159626 307727 159629
rect 307661 159624 310040 159626
rect 307661 159568 307666 159624
rect 307722 159568 310040 159624
rect 307661 159566 310040 159568
rect 307661 159563 307727 159566
rect 214649 159490 214715 159493
rect 214649 159488 217242 159490
rect 214649 159432 214654 159488
rect 214710 159432 217242 159488
rect 214649 159430 217242 159432
rect 214649 159427 214715 159430
rect 217182 159052 217242 159430
rect 324313 159354 324379 159357
rect 321908 159352 324379 159354
rect 321908 159296 324318 159352
rect 324374 159296 324379 159352
rect 321908 159294 324379 159296
rect 324313 159291 324379 159294
rect 252001 159218 252067 159221
rect 248952 159216 252067 159218
rect 248952 159160 252006 159216
rect 252062 159160 252067 159216
rect 248952 159158 252067 159160
rect 252001 159155 252067 159158
rect 306557 159082 306623 159085
rect 306557 159080 310040 159082
rect 306557 159024 306562 159080
rect 306618 159024 310040 159080
rect 306557 159022 310040 159024
rect 306557 159019 306623 159022
rect 251173 158810 251239 158813
rect 248952 158808 251239 158810
rect 248952 158752 251178 158808
rect 251234 158752 251239 158808
rect 248952 158750 251239 158752
rect 251173 158747 251239 158750
rect 213913 158674 213979 158677
rect 307569 158674 307635 158677
rect 213913 158672 217242 158674
rect 213913 158616 213918 158672
rect 213974 158616 217242 158672
rect 213913 158614 217242 158616
rect 213913 158611 213979 158614
rect 217182 158372 217242 158614
rect 307569 158672 310040 158674
rect 307569 158616 307574 158672
rect 307630 158616 310040 158672
rect 307569 158614 310040 158616
rect 307569 158611 307635 158614
rect 324313 158538 324379 158541
rect 321908 158536 324379 158538
rect 321908 158480 324318 158536
rect 324374 158480 324379 158536
rect 321908 158478 324379 158480
rect 324313 158475 324379 158478
rect 249885 158266 249951 158269
rect 248952 158264 249951 158266
rect 248952 158208 249890 158264
rect 249946 158208 249951 158264
rect 248952 158206 249951 158208
rect 249885 158203 249951 158206
rect 306925 158266 306991 158269
rect 306925 158264 310040 158266
rect 306925 158208 306930 158264
rect 306986 158208 310040 158264
rect 306925 158206 310040 158208
rect 306925 158203 306991 158206
rect 214005 158130 214071 158133
rect 214005 158128 217242 158130
rect 214005 158072 214010 158128
rect 214066 158072 217242 158128
rect 214005 158070 217242 158072
rect 214005 158067 214071 158070
rect 217182 157692 217242 158070
rect 307661 157858 307727 157861
rect 324405 157858 324471 157861
rect 307661 157856 310040 157858
rect 248860 157754 249442 157814
rect 307661 157800 307666 157856
rect 307722 157800 310040 157856
rect 307661 157798 310040 157800
rect 321908 157856 324471 157858
rect 321908 157800 324410 157856
rect 324466 157800 324471 157856
rect 321908 157798 324471 157800
rect 307661 157795 307727 157798
rect 324405 157795 324471 157798
rect 249382 157450 249442 157754
rect 269062 157450 269068 157452
rect 249382 157390 269068 157450
rect 269062 157388 269068 157390
rect 269132 157388 269138 157452
rect 305729 157450 305795 157453
rect 305729 157448 310040 157450
rect 305729 157392 305734 157448
rect 305790 157392 310040 157448
rect 305729 157390 310040 157392
rect 305729 157387 305795 157390
rect 213913 157314 213979 157317
rect 252461 157314 252527 157317
rect 213913 157312 217242 157314
rect 213913 157256 213918 157312
rect 213974 157256 217242 157312
rect 213913 157254 217242 157256
rect 248952 157312 252527 157314
rect 248952 157256 252466 157312
rect 252522 157256 252527 157312
rect 248952 157254 252527 157256
rect 213913 157251 213979 157254
rect 217182 157148 217242 157254
rect 252461 157251 252527 157254
rect 307477 157042 307543 157045
rect 322933 157042 322999 157045
rect 307477 157040 310040 157042
rect 307477 156984 307482 157040
rect 307538 156984 310040 157040
rect 307477 156982 310040 156984
rect 321908 157040 322999 157042
rect 321908 156984 322938 157040
rect 322994 156984 322999 157040
rect 321908 156982 322999 156984
rect 307477 156979 307543 156982
rect 322933 156979 322999 156982
rect 214005 156906 214071 156909
rect 252461 156906 252527 156909
rect 214005 156904 217242 156906
rect 214005 156848 214010 156904
rect 214066 156848 217242 156904
rect 214005 156846 217242 156848
rect 248952 156904 252527 156906
rect 248952 156848 252466 156904
rect 252522 156848 252527 156904
rect 248952 156846 252527 156848
rect 214005 156843 214071 156846
rect 217182 156468 217242 156846
rect 252461 156843 252527 156846
rect 307569 156634 307635 156637
rect 307569 156632 310040 156634
rect 307569 156576 307574 156632
rect 307630 156576 310040 156632
rect 307569 156574 310040 156576
rect 307569 156571 307635 156574
rect 252369 156362 252435 156365
rect 324313 156362 324379 156365
rect 248952 156360 252435 156362
rect 248952 156304 252374 156360
rect 252430 156304 252435 156360
rect 248952 156302 252435 156304
rect 321908 156360 324379 156362
rect 321908 156304 324318 156360
rect 324374 156304 324379 156360
rect 321908 156302 324379 156304
rect 252369 156299 252435 156302
rect 324313 156299 324379 156302
rect 307661 156226 307727 156229
rect 307661 156224 310040 156226
rect 307661 156168 307666 156224
rect 307722 156168 310040 156224
rect 307661 156166 310040 156168
rect 307661 156163 307727 156166
rect 252461 155954 252527 155957
rect 248952 155952 252527 155954
rect 248952 155896 252466 155952
rect 252522 155896 252527 155952
rect 248952 155894 252527 155896
rect 252461 155891 252527 155894
rect 213913 155546 213979 155549
rect 213913 155544 217242 155546
rect 213913 155488 213918 155544
rect 213974 155488 217242 155544
rect 213913 155486 217242 155488
rect 213913 155483 213979 155486
rect 217182 155108 217242 155486
rect 217366 155413 217426 155788
rect 307293 155682 307359 155685
rect 307293 155680 310040 155682
rect 307293 155624 307298 155680
rect 307354 155624 310040 155680
rect 307293 155622 310040 155624
rect 307293 155619 307359 155622
rect 324313 155546 324379 155549
rect 321908 155544 324379 155546
rect 321908 155488 324318 155544
rect 324374 155488 324379 155544
rect 321908 155486 324379 155488
rect 324313 155483 324379 155486
rect 217317 155408 217426 155413
rect 251449 155410 251515 155413
rect 217317 155352 217322 155408
rect 217378 155352 217426 155408
rect 217317 155350 217426 155352
rect 248952 155408 251515 155410
rect 248952 155352 251454 155408
rect 251510 155352 251515 155408
rect 248952 155350 251515 155352
rect 217317 155347 217383 155350
rect 251449 155347 251515 155350
rect 250437 155274 250503 155277
rect 258390 155274 258396 155276
rect 250437 155272 258396 155274
rect 250437 155216 250442 155272
rect 250498 155216 258396 155272
rect 250437 155214 258396 155216
rect 250437 155211 250503 155214
rect 258390 155212 258396 155214
rect 258460 155212 258466 155276
rect 307661 155274 307727 155277
rect 307661 155272 310040 155274
rect 307661 155216 307666 155272
rect 307722 155216 310040 155272
rect 307661 155214 310040 155216
rect 307661 155211 307727 155214
rect 252369 155002 252435 155005
rect 248952 155000 252435 155002
rect 248952 154944 252374 155000
rect 252430 154944 252435 155000
rect 248952 154942 252435 154944
rect 252369 154939 252435 154942
rect 306557 154866 306623 154869
rect 306557 154864 310040 154866
rect 306557 154808 306562 154864
rect 306618 154808 310040 154864
rect 306557 154806 310040 154808
rect 306557 154803 306623 154806
rect 217317 154730 217383 154733
rect 324405 154730 324471 154733
rect 200070 154728 217383 154730
rect 200070 154672 217322 154728
rect 217378 154672 217383 154728
rect 200070 154670 217383 154672
rect 321908 154728 324471 154730
rect 321908 154672 324410 154728
rect 324466 154672 324471 154728
rect 321908 154670 324471 154672
rect 166206 154532 166212 154596
rect 166276 154594 166282 154596
rect 200070 154594 200130 154670
rect 217317 154667 217383 154670
rect 324405 154667 324471 154670
rect 166276 154534 200130 154594
rect 166276 154532 166282 154534
rect 252461 154458 252527 154461
rect 248952 154456 252527 154458
rect 214005 153914 214071 153917
rect 217182 153914 217242 154428
rect 248952 154400 252466 154456
rect 252522 154400 252527 154456
rect 248952 154398 252527 154400
rect 252461 154395 252527 154398
rect 306557 154458 306623 154461
rect 306557 154456 310040 154458
rect 306557 154400 306562 154456
rect 306618 154400 310040 154456
rect 306557 154398 310040 154400
rect 306557 154395 306623 154398
rect 252369 154050 252435 154053
rect 324313 154050 324379 154053
rect 248952 154048 252435 154050
rect 248952 153992 252374 154048
rect 252430 153992 252435 154048
rect 321908 154048 324379 154050
rect 248952 153990 252435 153992
rect 252369 153987 252435 153990
rect 309550 153946 310132 154006
rect 321908 153992 324318 154048
rect 324374 153992 324379 154048
rect 321908 153990 324379 153992
rect 324313 153987 324379 153990
rect 309550 153914 309610 153946
rect 214005 153912 217242 153914
rect 214005 153856 214010 153912
rect 214066 153856 217242 153912
rect 214005 153854 217242 153856
rect 296670 153854 309610 153914
rect 214005 153851 214071 153854
rect 213913 153506 213979 153509
rect 217182 153506 217242 153748
rect 213913 153504 217242 153506
rect 213913 153448 213918 153504
rect 213974 153448 217242 153504
rect 213913 153446 217242 153448
rect 213913 153443 213979 153446
rect 248860 153402 249442 153462
rect 258574 153444 258580 153508
rect 258644 153506 258650 153508
rect 296670 153506 296730 153854
rect 307661 153642 307727 153645
rect 307661 153640 310040 153642
rect 307661 153584 307666 153640
rect 307722 153584 310040 153640
rect 307661 153582 310040 153584
rect 307661 153579 307727 153582
rect 258644 153446 296730 153506
rect 258644 153444 258650 153446
rect 249382 153370 249442 153402
rect 266302 153370 266308 153372
rect 249382 153310 266308 153370
rect 266302 153308 266308 153310
rect 266372 153308 266378 153372
rect 306649 153234 306715 153237
rect 324313 153234 324379 153237
rect 306649 153232 310040 153234
rect 306649 153176 306654 153232
rect 306710 153176 310040 153232
rect 306649 153174 310040 153176
rect 321908 153232 324379 153234
rect 321908 153176 324318 153232
rect 324374 153176 324379 153232
rect 321908 153174 324379 153176
rect 306649 153171 306715 153174
rect 324313 153171 324379 153174
rect 252461 153098 252527 153101
rect 248952 153096 252527 153098
rect 213177 152690 213243 152693
rect 217182 152690 217242 153068
rect 248952 153040 252466 153096
rect 252522 153040 252527 153096
rect 248952 153038 252527 153040
rect 252461 153035 252527 153038
rect 252553 152690 252619 152693
rect 213177 152688 217242 152690
rect 213177 152632 213182 152688
rect 213238 152632 217242 152688
rect 213177 152630 217242 152632
rect 248952 152688 252619 152690
rect 248952 152632 252558 152688
rect 252614 152632 252619 152688
rect 248952 152630 252619 152632
rect 213177 152627 213243 152630
rect 252553 152627 252619 152630
rect 307477 152690 307543 152693
rect 579797 152690 579863 152693
rect 583520 152690 584960 152780
rect 307477 152688 310040 152690
rect 307477 152632 307482 152688
rect 307538 152632 310040 152688
rect 307477 152630 310040 152632
rect 579797 152688 584960 152690
rect 579797 152632 579802 152688
rect 579858 152632 584960 152688
rect 579797 152630 584960 152632
rect 307477 152627 307543 152630
rect 579797 152627 579863 152630
rect 583520 152540 584960 152630
rect 214373 152146 214439 152149
rect 217182 152146 217242 152524
rect 324405 152418 324471 152421
rect 321908 152416 324471 152418
rect 321908 152360 324410 152416
rect 324466 152360 324471 152416
rect 321908 152358 324471 152360
rect 324405 152355 324471 152358
rect 307569 152282 307635 152285
rect 307569 152280 310040 152282
rect 307569 152224 307574 152280
rect 307630 152224 310040 152280
rect 307569 152222 310040 152224
rect 307569 152219 307635 152222
rect 252277 152146 252343 152149
rect 214373 152144 217242 152146
rect 214373 152088 214378 152144
rect 214434 152088 217242 152144
rect 214373 152086 217242 152088
rect 248952 152144 252343 152146
rect 248952 152088 252282 152144
rect 252338 152088 252343 152144
rect 248952 152086 252343 152088
rect 214373 152083 214439 152086
rect 252277 152083 252343 152086
rect 213913 152010 213979 152013
rect 213913 152008 217242 152010
rect 213913 151952 213918 152008
rect 213974 151952 217242 152008
rect 213913 151950 217242 151952
rect 213913 151947 213979 151950
rect 217182 151844 217242 151950
rect 307661 151874 307727 151877
rect 307661 151872 310040 151874
rect 307661 151816 307666 151872
rect 307722 151816 310040 151872
rect 307661 151814 310040 151816
rect 307661 151811 307727 151814
rect 252461 151738 252527 151741
rect 324313 151738 324379 151741
rect 248952 151736 252527 151738
rect 248952 151680 252466 151736
rect 252522 151680 252527 151736
rect 248952 151678 252527 151680
rect 321908 151736 324379 151738
rect 321908 151680 324318 151736
rect 324374 151680 324379 151736
rect 321908 151678 324379 151680
rect 252461 151675 252527 151678
rect 324313 151675 324379 151678
rect 307293 151466 307359 151469
rect 307293 151464 310040 151466
rect 307293 151408 307298 151464
rect 307354 151408 310040 151464
rect 307293 151406 310040 151408
rect 307293 151403 307359 151406
rect 252001 151194 252067 151197
rect 248952 151192 252067 151194
rect 214005 150922 214071 150925
rect 217182 150922 217242 151164
rect 248952 151136 252006 151192
rect 252062 151136 252067 151192
rect 248952 151134 252067 151136
rect 252001 151131 252067 151134
rect 306925 151058 306991 151061
rect 306925 151056 310040 151058
rect 306925 151000 306930 151056
rect 306986 151000 310040 151056
rect 306925 150998 310040 151000
rect 306925 150995 306991 150998
rect 325877 150922 325943 150925
rect 214005 150920 217242 150922
rect 214005 150864 214010 150920
rect 214066 150864 217242 150920
rect 214005 150862 217242 150864
rect 321908 150920 325943 150922
rect 321908 150864 325882 150920
rect 325938 150864 325943 150920
rect 321908 150862 325943 150864
rect 214005 150859 214071 150862
rect 325877 150859 325943 150862
rect 214649 150786 214715 150789
rect 249793 150786 249859 150789
rect 214649 150784 217426 150786
rect 214649 150728 214654 150784
rect 214710 150728 217426 150784
rect 214649 150726 217426 150728
rect 248952 150784 249859 150786
rect 248952 150728 249798 150784
rect 249854 150728 249859 150784
rect 248952 150726 249859 150728
rect 214649 150723 214715 150726
rect 217366 150484 217426 150726
rect 249793 150723 249859 150726
rect 307661 150650 307727 150653
rect 307661 150648 310040 150650
rect 307661 150592 307666 150648
rect 307722 150592 310040 150648
rect 307661 150590 310040 150592
rect 307661 150587 307727 150590
rect 252277 150242 252343 150245
rect 248952 150240 252343 150242
rect 248952 150184 252282 150240
rect 252338 150184 252343 150240
rect 248952 150182 252343 150184
rect 252277 150179 252343 150182
rect 307661 150242 307727 150245
rect 307661 150240 310040 150242
rect 307661 150184 307666 150240
rect 307722 150184 310040 150240
rect 307661 150182 310040 150184
rect 307661 150179 307727 150182
rect 213913 150106 213979 150109
rect 324313 150106 324379 150109
rect 213913 150104 217242 150106
rect 213913 150048 213918 150104
rect 213974 150048 217242 150104
rect 213913 150046 217242 150048
rect 321908 150104 324379 150106
rect 321908 150048 324318 150104
rect 324374 150048 324379 150104
rect 321908 150046 324379 150048
rect 213913 150043 213979 150046
rect -960 149834 480 149924
rect 3509 149834 3575 149837
rect -960 149832 3575 149834
rect -960 149776 3514 149832
rect 3570 149776 3575 149832
rect 217182 149804 217242 150046
rect 324313 150043 324379 150046
rect 252461 149834 252527 149837
rect 248952 149832 252527 149834
rect -960 149774 3575 149776
rect 248952 149776 252466 149832
rect 252522 149776 252527 149832
rect 248952 149774 252527 149776
rect -960 149684 480 149774
rect 3509 149771 3575 149774
rect 252461 149771 252527 149774
rect 307385 149834 307451 149837
rect 307385 149832 310040 149834
rect 307385 149776 307390 149832
rect 307446 149776 310040 149832
rect 307385 149774 310040 149776
rect 307385 149771 307451 149774
rect 214557 149562 214623 149565
rect 214557 149560 217242 149562
rect 214557 149504 214562 149560
rect 214618 149504 217242 149560
rect 214557 149502 217242 149504
rect 214557 149499 214623 149502
rect 217182 149124 217242 149502
rect 324405 149426 324471 149429
rect 321908 149424 324471 149426
rect 321908 149368 324410 149424
rect 324466 149368 324471 149424
rect 321908 149366 324471 149368
rect 324405 149363 324471 149366
rect 252369 149290 252435 149293
rect 248952 149288 252435 149290
rect 248952 149232 252374 149288
rect 252430 149232 252435 149288
rect 248952 149230 252435 149232
rect 252369 149227 252435 149230
rect 307569 149290 307635 149293
rect 307569 149288 310040 149290
rect 307569 149232 307574 149288
rect 307630 149232 310040 149288
rect 307569 149230 310040 149232
rect 307569 149227 307635 149230
rect 252829 148882 252895 148885
rect 248952 148880 252895 148882
rect 248952 148824 252834 148880
rect 252890 148824 252895 148880
rect 248952 148822 252895 148824
rect 252829 148819 252895 148822
rect 306557 148882 306623 148885
rect 306557 148880 310040 148882
rect 306557 148824 306562 148880
rect 306618 148824 310040 148880
rect 306557 148822 310040 148824
rect 306557 148819 306623 148822
rect 213913 148746 213979 148749
rect 213913 148744 217242 148746
rect 213913 148688 213918 148744
rect 213974 148688 217242 148744
rect 213913 148686 217242 148688
rect 213913 148683 213979 148686
rect 217182 148444 217242 148686
rect 324313 148610 324379 148613
rect 321908 148608 324379 148610
rect 321908 148552 324318 148608
rect 324374 148552 324379 148608
rect 321908 148550 324379 148552
rect 324313 148547 324379 148550
rect 307661 148474 307727 148477
rect 307661 148472 310040 148474
rect 307661 148416 307666 148472
rect 307722 148416 310040 148472
rect 307661 148414 310040 148416
rect 307661 148411 307727 148414
rect 252461 148338 252527 148341
rect 303521 148338 303587 148341
rect 321737 148338 321803 148341
rect 248952 148336 252527 148338
rect 248952 148280 252466 148336
rect 252522 148280 252527 148336
rect 248952 148278 252527 148280
rect 252461 148275 252527 148278
rect 258030 148336 303587 148338
rect 258030 148280 303526 148336
rect 303582 148280 303587 148336
rect 258030 148278 303587 148280
rect 251766 148140 251772 148204
rect 251836 148202 251842 148204
rect 258030 148202 258090 148278
rect 303521 148275 303587 148278
rect 321694 148336 321803 148338
rect 321694 148280 321742 148336
rect 321798 148280 321803 148336
rect 321694 148275 321803 148280
rect 251836 148142 258090 148202
rect 251836 148140 251842 148142
rect 213913 148066 213979 148069
rect 213913 148064 217242 148066
rect 213913 148008 213918 148064
rect 213974 148008 217242 148064
rect 213913 148006 217242 148008
rect 213913 148003 213979 148006
rect 217182 147900 217242 148006
rect 309550 147962 310132 148022
rect 252369 147930 252435 147933
rect 248952 147928 252435 147930
rect 248952 147872 252374 147928
rect 252430 147872 252435 147928
rect 248952 147870 252435 147872
rect 252369 147867 252435 147870
rect 305913 147930 305979 147933
rect 309550 147930 309610 147962
rect 305913 147928 309610 147930
rect 305913 147872 305918 147928
rect 305974 147872 309610 147928
rect 305913 147870 309610 147872
rect 305913 147867 305979 147870
rect 321694 147764 321754 148275
rect 307477 147658 307543 147661
rect 307477 147656 310040 147658
rect 307477 147600 307482 147656
rect 307538 147600 310040 147656
rect 307477 147598 310040 147600
rect 307477 147595 307543 147598
rect 255262 147522 255268 147524
rect 248952 147462 255268 147522
rect 255262 147460 255268 147462
rect 255332 147460 255338 147524
rect 307293 147250 307359 147253
rect 307293 147248 310040 147250
rect 214005 146706 214071 146709
rect 217182 146706 217242 147220
rect 307293 147192 307298 147248
rect 307354 147192 310040 147248
rect 307293 147190 310040 147192
rect 307293 147187 307359 147190
rect 324313 147114 324379 147117
rect 321908 147112 324379 147114
rect 321908 147056 324318 147112
rect 324374 147056 324379 147112
rect 321908 147054 324379 147056
rect 324313 147051 324379 147054
rect 251265 146978 251331 146981
rect 248952 146976 251331 146978
rect 248952 146920 251270 146976
rect 251326 146920 251331 146976
rect 248952 146918 251331 146920
rect 251265 146915 251331 146918
rect 306925 146842 306991 146845
rect 306925 146840 310040 146842
rect 306925 146784 306930 146840
rect 306986 146784 310040 146840
rect 306925 146782 310040 146784
rect 306925 146779 306991 146782
rect 214005 146704 217242 146706
rect 214005 146648 214010 146704
rect 214066 146648 217242 146704
rect 214005 146646 217242 146648
rect 214005 146643 214071 146646
rect 252461 146570 252527 146573
rect 248952 146568 252527 146570
rect 213913 146434 213979 146437
rect 213913 146432 216874 146434
rect 213913 146376 213918 146432
rect 213974 146376 216874 146432
rect 213913 146374 216874 146376
rect 213913 146371 213979 146374
rect 216814 146298 216874 146374
rect 217366 146298 217426 146540
rect 248952 146512 252466 146568
rect 252522 146512 252527 146568
rect 248952 146510 252527 146512
rect 252461 146507 252527 146510
rect 307702 146372 307708 146436
rect 307772 146434 307778 146436
rect 307772 146374 310040 146434
rect 307772 146372 307778 146374
rect 216814 146238 217426 146298
rect 252185 146298 252251 146301
rect 258390 146298 258396 146300
rect 252185 146296 258396 146298
rect 252185 146240 252190 146296
rect 252246 146240 258396 146296
rect 252185 146238 258396 146240
rect 252185 146235 252251 146238
rect 258390 146236 258396 146238
rect 258460 146236 258466 146300
rect 324313 146298 324379 146301
rect 321908 146296 324379 146298
rect 321908 146240 324318 146296
rect 324374 146240 324379 146296
rect 321908 146238 324379 146240
rect 324313 146235 324379 146238
rect 252461 146026 252527 146029
rect 248952 146024 252527 146026
rect 248952 145968 252466 146024
rect 252522 145968 252527 146024
rect 248952 145966 252527 145968
rect 252461 145963 252527 145966
rect 307109 145890 307175 145893
rect 307109 145888 310040 145890
rect 214005 145346 214071 145349
rect 217182 145346 217242 145860
rect 307109 145832 307114 145888
rect 307170 145832 310040 145888
rect 307109 145830 310040 145832
rect 307109 145827 307175 145830
rect 252369 145618 252435 145621
rect 248952 145616 252435 145618
rect 248952 145560 252374 145616
rect 252430 145560 252435 145616
rect 248952 145558 252435 145560
rect 252369 145555 252435 145558
rect 265617 145618 265683 145621
rect 307702 145618 307708 145620
rect 265617 145616 307708 145618
rect 265617 145560 265622 145616
rect 265678 145560 307708 145616
rect 265617 145558 307708 145560
rect 265617 145555 265683 145558
rect 307702 145556 307708 145558
rect 307772 145556 307778 145620
rect 324405 145482 324471 145485
rect 321908 145480 324471 145482
rect 214005 145344 217242 145346
rect 214005 145288 214010 145344
rect 214066 145288 217242 145344
rect 214005 145286 217242 145288
rect 309550 145378 310132 145438
rect 321908 145424 324410 145480
rect 324466 145424 324471 145480
rect 321908 145422 324471 145424
rect 324405 145419 324471 145422
rect 214005 145283 214071 145286
rect 213913 144938 213979 144941
rect 217366 144938 217426 145180
rect 252277 145074 252343 145077
rect 248952 145072 252343 145074
rect 248952 145016 252282 145072
rect 252338 145016 252343 145072
rect 248952 145014 252343 145016
rect 252277 145011 252343 145014
rect 305637 145074 305703 145077
rect 309550 145074 309610 145378
rect 305637 145072 309610 145074
rect 305637 145016 305642 145072
rect 305698 145016 309610 145072
rect 305637 145014 309610 145016
rect 305637 145011 305703 145014
rect 309734 144970 310132 145030
rect 213913 144936 217426 144938
rect 213913 144880 213918 144936
rect 213974 144880 217426 144936
rect 213913 144878 217426 144880
rect 307385 144938 307451 144941
rect 309734 144938 309794 144970
rect 307385 144936 309794 144938
rect 307385 144880 307390 144936
rect 307446 144880 309794 144936
rect 307385 144878 309794 144880
rect 213913 144875 213979 144878
rect 307385 144875 307451 144878
rect 324313 144802 324379 144805
rect 321908 144800 324379 144802
rect 321908 144744 324318 144800
rect 324374 144744 324379 144800
rect 321908 144742 324379 144744
rect 324313 144739 324379 144742
rect 307477 144666 307543 144669
rect 307477 144664 310040 144666
rect 248860 144562 249442 144622
rect 307477 144608 307482 144664
rect 307538 144608 310040 144664
rect 307477 144606 310040 144608
rect 307477 144603 307543 144606
rect 249382 144530 249442 144562
rect 263542 144530 263548 144532
rect 214005 143986 214071 143989
rect 217182 143986 217242 144500
rect 249382 144470 263548 144530
rect 263542 144468 263548 144470
rect 263612 144468 263618 144532
rect 307569 144258 307635 144261
rect 307569 144256 310040 144258
rect 307569 144200 307574 144256
rect 307630 144200 310040 144256
rect 307569 144198 310040 144200
rect 307569 144195 307635 144198
rect 252461 144122 252527 144125
rect 248952 144120 252527 144122
rect 248952 144064 252466 144120
rect 252522 144064 252527 144120
rect 248952 144062 252527 144064
rect 252461 144059 252527 144062
rect 324405 143986 324471 143989
rect 214005 143984 217242 143986
rect 214005 143928 214010 143984
rect 214066 143928 217242 143984
rect 214005 143926 217242 143928
rect 321908 143984 324471 143986
rect 321908 143928 324410 143984
rect 324466 143928 324471 143984
rect 321908 143926 324471 143928
rect 214005 143923 214071 143926
rect 324405 143923 324471 143926
rect 307661 143850 307727 143853
rect 307661 143848 310040 143850
rect 213913 143578 213979 143581
rect 217366 143578 217426 143820
rect 307661 143792 307666 143848
rect 307722 143792 310040 143848
rect 307661 143790 310040 143792
rect 307661 143787 307727 143790
rect 250437 143714 250503 143717
rect 248952 143712 250503 143714
rect 248952 143656 250442 143712
rect 250498 143656 250503 143712
rect 248952 143654 250503 143656
rect 250437 143651 250503 143654
rect 213913 143576 217426 143578
rect 213913 143520 213918 143576
rect 213974 143520 217426 143576
rect 213913 143518 217426 143520
rect 213913 143515 213979 143518
rect 306557 143442 306623 143445
rect 306557 143440 310040 143442
rect 306557 143384 306562 143440
rect 306618 143384 310040 143440
rect 306557 143382 310040 143384
rect 306557 143379 306623 143382
rect 217182 142762 217242 143276
rect 252461 143170 252527 143173
rect 324313 143170 324379 143173
rect 248952 143168 252527 143170
rect 248952 143112 252466 143168
rect 252522 143112 252527 143168
rect 248952 143110 252527 143112
rect 321908 143168 324379 143170
rect 321908 143112 324318 143168
rect 324374 143112 324379 143168
rect 321908 143110 324379 143112
rect 252461 143107 252527 143110
rect 324313 143107 324379 143110
rect 307569 143034 307635 143037
rect 307569 143032 310040 143034
rect 307569 142976 307574 143032
rect 307630 142976 310040 143032
rect 307569 142974 310040 142976
rect 307569 142971 307635 142974
rect 252185 142762 252251 142765
rect 200070 142702 217242 142762
rect 248952 142760 252251 142762
rect 248952 142704 252190 142760
rect 252246 142704 252251 142760
rect 248952 142702 252251 142704
rect 168966 142156 168972 142220
rect 169036 142218 169042 142220
rect 200070 142218 200130 142702
rect 252185 142699 252251 142702
rect 169036 142158 200130 142218
rect 213913 142218 213979 142221
rect 217182 142218 217242 142596
rect 307661 142490 307727 142493
rect 324405 142490 324471 142493
rect 307661 142488 310040 142490
rect 307661 142432 307666 142488
rect 307722 142432 310040 142488
rect 307661 142430 310040 142432
rect 321908 142488 324471 142490
rect 321908 142432 324410 142488
rect 324466 142432 324471 142488
rect 321908 142430 324471 142432
rect 307661 142427 307727 142430
rect 324405 142427 324471 142430
rect 251950 142292 251956 142356
rect 252020 142354 252026 142356
rect 258993 142354 259059 142357
rect 252020 142352 259059 142354
rect 252020 142296 258998 142352
rect 259054 142296 259059 142352
rect 252020 142294 259059 142296
rect 252020 142292 252026 142294
rect 258993 142291 259059 142294
rect 252369 142218 252435 142221
rect 213913 142216 217242 142218
rect 213913 142160 213918 142216
rect 213974 142160 217242 142216
rect 213913 142158 217242 142160
rect 248952 142216 252435 142218
rect 248952 142160 252374 142216
rect 252430 142160 252435 142216
rect 248952 142158 252435 142160
rect 169036 142156 169042 142158
rect 213913 142155 213979 142158
rect 252369 142155 252435 142158
rect 306557 142082 306623 142085
rect 306557 142080 310040 142082
rect 306557 142024 306562 142080
rect 306618 142024 310040 142080
rect 306557 142022 310040 142024
rect 306557 142019 306623 142022
rect 214005 141402 214071 141405
rect 217182 141402 217242 141916
rect 248860 141706 249442 141766
rect 249382 141674 249442 141706
rect 307569 141674 307635 141677
rect 324313 141674 324379 141677
rect 249382 141614 258090 141674
rect 252461 141402 252527 141405
rect 214005 141400 217242 141402
rect 214005 141344 214010 141400
rect 214066 141344 217242 141400
rect 214005 141342 217242 141344
rect 248952 141400 252527 141402
rect 248952 141344 252466 141400
rect 252522 141344 252527 141400
rect 248952 141342 252527 141344
rect 214005 141339 214071 141342
rect 252461 141339 252527 141342
rect 213913 140994 213979 140997
rect 217182 140994 217242 141236
rect 213913 140992 217242 140994
rect 213913 140936 213918 140992
rect 213974 140936 217242 140992
rect 213913 140934 217242 140936
rect 213913 140931 213979 140934
rect 251357 140858 251423 140861
rect 248952 140856 251423 140858
rect 248952 140800 251362 140856
rect 251418 140800 251423 140856
rect 248952 140798 251423 140800
rect 258030 140858 258090 141614
rect 307569 141672 310040 141674
rect 307569 141616 307574 141672
rect 307630 141616 310040 141672
rect 307569 141614 310040 141616
rect 321908 141672 324379 141674
rect 321908 141616 324318 141672
rect 324374 141616 324379 141672
rect 321908 141614 324379 141616
rect 307569 141611 307635 141614
rect 324313 141611 324379 141614
rect 307661 141266 307727 141269
rect 307661 141264 310040 141266
rect 307661 141208 307666 141264
rect 307722 141208 310040 141264
rect 307661 141206 310040 141208
rect 307661 141203 307727 141206
rect 267774 140858 267780 140860
rect 258030 140798 267780 140858
rect 251357 140795 251423 140798
rect 267774 140796 267780 140798
rect 267844 140796 267850 140860
rect 306741 140858 306807 140861
rect 324405 140858 324471 140861
rect 306741 140856 310040 140858
rect 306741 140800 306746 140856
rect 306802 140800 310040 140856
rect 306741 140798 310040 140800
rect 321908 140856 324471 140858
rect 321908 140800 324410 140856
rect 324466 140800 324471 140856
rect 321908 140798 324471 140800
rect 306741 140795 306807 140798
rect 324405 140795 324471 140798
rect 214005 140042 214071 140045
rect 217182 140042 217242 140556
rect 256734 140450 256740 140452
rect 248952 140390 256740 140450
rect 256734 140388 256740 140390
rect 256804 140388 256810 140452
rect 307201 140450 307267 140453
rect 307201 140448 310040 140450
rect 307201 140392 307206 140448
rect 307262 140392 310040 140448
rect 307201 140390 310040 140392
rect 307201 140387 307267 140390
rect 324313 140178 324379 140181
rect 321908 140176 324379 140178
rect 321908 140120 324318 140176
rect 324374 140120 324379 140176
rect 321908 140118 324379 140120
rect 324313 140115 324379 140118
rect 214005 140040 217242 140042
rect 214005 139984 214010 140040
rect 214066 139984 217242 140040
rect 214005 139982 217242 139984
rect 306925 140042 306991 140045
rect 306925 140040 310040 140042
rect 306925 139984 306930 140040
rect 306986 139984 310040 140040
rect 306925 139982 310040 139984
rect 214005 139979 214071 139982
rect 306925 139979 306991 139982
rect 252461 139906 252527 139909
rect 248952 139904 252527 139906
rect 213913 139634 213979 139637
rect 217182 139634 217242 139876
rect 248952 139848 252466 139904
rect 252522 139848 252527 139904
rect 248952 139846 252527 139848
rect 252461 139843 252527 139846
rect 213913 139632 217242 139634
rect 213913 139576 213918 139632
rect 213974 139576 217242 139632
rect 213913 139574 217242 139576
rect 307293 139634 307359 139637
rect 307293 139632 310040 139634
rect 307293 139576 307298 139632
rect 307354 139576 310040 139632
rect 307293 139574 310040 139576
rect 213913 139571 213979 139574
rect 307293 139571 307359 139574
rect 252369 139498 252435 139501
rect 248952 139496 252435 139498
rect 248952 139440 252374 139496
rect 252430 139440 252435 139496
rect 248952 139438 252435 139440
rect 252369 139435 252435 139438
rect 324313 139362 324379 139365
rect 583520 139362 584960 139452
rect 321908 139360 324379 139362
rect 321908 139304 324318 139360
rect 324374 139304 324379 139360
rect 321908 139302 324379 139304
rect 324313 139299 324379 139302
rect 583342 139302 584960 139362
rect 583342 139226 583402 139302
rect 583520 139226 584960 139302
rect 583342 139212 584960 139226
rect 214465 138818 214531 138821
rect 217182 138818 217242 139196
rect 583342 139166 583586 139212
rect 306557 139090 306623 139093
rect 306557 139088 310040 139090
rect 306557 139032 306562 139088
rect 306618 139032 310040 139088
rect 306557 139030 310040 139032
rect 306557 139027 306623 139030
rect 248860 138850 249442 138910
rect 214465 138816 217242 138818
rect 214465 138760 214470 138816
rect 214526 138760 217242 138816
rect 214465 138758 217242 138760
rect 249382 138818 249442 138850
rect 263726 138818 263732 138820
rect 249382 138758 263732 138818
rect 214465 138755 214531 138758
rect 263726 138756 263732 138758
rect 263796 138756 263802 138820
rect 307569 138682 307635 138685
rect 307569 138680 310040 138682
rect 213913 138138 213979 138141
rect 217182 138138 217242 138652
rect 307569 138624 307574 138680
rect 307630 138624 310040 138680
rect 307569 138622 310040 138624
rect 307569 138619 307635 138622
rect 252277 138546 252343 138549
rect 324405 138546 324471 138549
rect 248952 138544 252343 138546
rect 248952 138488 252282 138544
rect 252338 138488 252343 138544
rect 248952 138486 252343 138488
rect 321908 138544 324471 138546
rect 321908 138488 324410 138544
rect 324466 138488 324471 138544
rect 321908 138486 324471 138488
rect 252277 138483 252343 138486
rect 324405 138483 324471 138486
rect 307661 138274 307727 138277
rect 307661 138272 310040 138274
rect 307661 138216 307666 138272
rect 307722 138216 310040 138272
rect 307661 138214 310040 138216
rect 307661 138211 307727 138214
rect 213913 138136 217242 138138
rect 213913 138080 213918 138136
rect 213974 138080 217242 138136
rect 213913 138078 217242 138080
rect 213913 138075 213979 138078
rect 342110 138076 342116 138140
rect 342180 138138 342186 138140
rect 583526 138138 583586 139166
rect 342180 138078 583586 138138
rect 342180 138076 342186 138078
rect 252369 138002 252435 138005
rect 248952 138000 252435 138002
rect 214649 137458 214715 137461
rect 217182 137458 217242 137972
rect 248952 137944 252374 138000
rect 252430 137944 252435 138000
rect 248952 137942 252435 137944
rect 252369 137939 252435 137942
rect 307109 137866 307175 137869
rect 324313 137866 324379 137869
rect 307109 137864 310040 137866
rect 307109 137808 307114 137864
rect 307170 137808 310040 137864
rect 307109 137806 310040 137808
rect 321908 137864 324379 137866
rect 321908 137808 324318 137864
rect 324374 137808 324379 137864
rect 321908 137806 324379 137808
rect 307109 137803 307175 137806
rect 324313 137803 324379 137806
rect 252461 137594 252527 137597
rect 248952 137592 252527 137594
rect 248952 137536 252466 137592
rect 252522 137536 252527 137592
rect 248952 137534 252527 137536
rect 252461 137531 252527 137534
rect 214649 137456 217242 137458
rect 214649 137400 214654 137456
rect 214710 137400 217242 137456
rect 214649 137398 217242 137400
rect 307569 137458 307635 137461
rect 307569 137456 310040 137458
rect 307569 137400 307574 137456
rect 307630 137400 310040 137456
rect 307569 137398 310040 137400
rect 214649 137395 214715 137398
rect 307569 137395 307635 137398
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 213913 136778 213979 136781
rect 217182 136778 217242 137292
rect 252277 137050 252343 137053
rect 248952 137048 252343 137050
rect 248952 136992 252282 137048
rect 252338 136992 252343 137048
rect 248952 136990 252343 136992
rect 252277 136987 252343 136990
rect 307661 137050 307727 137053
rect 324405 137050 324471 137053
rect 307661 137048 310040 137050
rect 307661 136992 307666 137048
rect 307722 136992 310040 137048
rect 307661 136990 310040 136992
rect 321908 137048 324471 137050
rect 321908 136992 324410 137048
rect 324466 136992 324471 137048
rect 321908 136990 324471 136992
rect 307661 136987 307727 136990
rect 324405 136987 324471 136990
rect 213913 136776 217242 136778
rect 213913 136720 213918 136776
rect 213974 136720 217242 136776
rect 213913 136718 217242 136720
rect 213913 136715 213979 136718
rect 252461 136642 252527 136645
rect 248952 136640 252527 136642
rect 217182 136098 217242 136612
rect 248952 136584 252466 136640
rect 252522 136584 252527 136640
rect 248952 136582 252527 136584
rect 252461 136579 252527 136582
rect 307477 136642 307543 136645
rect 307477 136640 310040 136642
rect 307477 136584 307482 136640
rect 307538 136584 310040 136640
rect 307477 136582 310040 136584
rect 307477 136579 307543 136582
rect 324313 136370 324379 136373
rect 321908 136368 324379 136370
rect 321908 136312 324318 136368
rect 324374 136312 324379 136368
rect 321908 136310 324379 136312
rect 324313 136307 324379 136310
rect 252001 136234 252067 136237
rect 248952 136232 252067 136234
rect 248952 136176 252006 136232
rect 252062 136176 252067 136232
rect 248952 136174 252067 136176
rect 252001 136171 252067 136174
rect 306557 136234 306623 136237
rect 306557 136232 310040 136234
rect 306557 136176 306562 136232
rect 306618 136176 310040 136232
rect 306557 136174 310040 136176
rect 306557 136171 306623 136174
rect 200070 136038 217242 136098
rect 166206 135492 166212 135556
rect 166276 135554 166282 135556
rect 200070 135554 200130 136038
rect 214005 135690 214071 135693
rect 217182 135690 217242 135932
rect 252277 135690 252343 135693
rect 214005 135688 217242 135690
rect 214005 135632 214010 135688
rect 214066 135632 217242 135688
rect 214005 135630 217242 135632
rect 248952 135688 252343 135690
rect 248952 135632 252282 135688
rect 252338 135632 252343 135688
rect 248952 135630 252343 135632
rect 214005 135627 214071 135630
rect 252277 135627 252343 135630
rect 307293 135690 307359 135693
rect 307293 135688 310040 135690
rect 307293 135632 307298 135688
rect 307354 135632 310040 135688
rect 307293 135630 310040 135632
rect 307293 135627 307359 135630
rect 166276 135494 200130 135554
rect 166276 135492 166282 135494
rect 213913 135418 213979 135421
rect 213913 135416 217242 135418
rect 213913 135360 213918 135416
rect 213974 135360 217242 135416
rect 213913 135358 217242 135360
rect 213913 135355 213979 135358
rect 217182 135252 217242 135358
rect 252369 135282 252435 135285
rect 248952 135280 252435 135282
rect 248952 135224 252374 135280
rect 252430 135224 252435 135280
rect 248952 135222 252435 135224
rect 252369 135219 252435 135222
rect 307661 135282 307727 135285
rect 321878 135282 321938 135524
rect 336774 135282 336780 135284
rect 307661 135280 310040 135282
rect 307661 135224 307666 135280
rect 307722 135224 310040 135280
rect 307661 135222 310040 135224
rect 321878 135222 336780 135282
rect 307661 135219 307727 135222
rect 336774 135220 336780 135222
rect 336844 135220 336850 135284
rect 307569 134874 307635 134877
rect 307569 134872 310040 134874
rect 307569 134816 307574 134872
rect 307630 134816 310040 134872
rect 307569 134814 310040 134816
rect 307569 134811 307635 134814
rect 252461 134738 252527 134741
rect 324313 134738 324379 134741
rect 248952 134736 252527 134738
rect 248952 134680 252466 134736
rect 252522 134680 252527 134736
rect 248952 134678 252527 134680
rect 321908 134736 324379 134738
rect 321908 134680 324318 134736
rect 324374 134680 324379 134736
rect 321908 134678 324379 134680
rect 252461 134675 252527 134678
rect 324313 134675 324379 134678
rect 214005 134330 214071 134333
rect 217182 134330 217242 134572
rect 307661 134466 307727 134469
rect 307661 134464 310040 134466
rect 307661 134408 307666 134464
rect 307722 134408 310040 134464
rect 307661 134406 310040 134408
rect 307661 134403 307727 134406
rect 252369 134330 252435 134333
rect 214005 134328 217242 134330
rect 214005 134272 214010 134328
rect 214066 134272 217242 134328
rect 214005 134270 217242 134272
rect 248952 134328 252435 134330
rect 248952 134272 252374 134328
rect 252430 134272 252435 134328
rect 248952 134270 252435 134272
rect 214005 134267 214071 134270
rect 252369 134267 252435 134270
rect 213913 134058 213979 134061
rect 213913 134056 217242 134058
rect 213913 134000 213918 134056
rect 213974 134000 217242 134056
rect 213913 133998 217242 134000
rect 213913 133995 213979 133998
rect 217182 133892 217242 133998
rect 302734 133996 302740 134060
rect 302804 134058 302810 134060
rect 325785 134058 325851 134061
rect 302804 133998 310040 134058
rect 321908 134056 325851 134058
rect 321908 134000 325790 134056
rect 325846 134000 325851 134056
rect 321908 133998 325851 134000
rect 302804 133996 302810 133998
rect 325785 133995 325851 133998
rect 252461 133786 252527 133789
rect 248952 133784 252527 133786
rect 248952 133728 252466 133784
rect 252522 133728 252527 133784
rect 248952 133726 252527 133728
rect 252461 133723 252527 133726
rect 307569 133650 307635 133653
rect 307569 133648 310040 133650
rect 307569 133592 307574 133648
rect 307630 133592 310040 133648
rect 307569 133590 310040 133592
rect 307569 133587 307635 133590
rect 252369 133378 252435 133381
rect 248952 133376 252435 133378
rect 214005 132834 214071 132837
rect 217182 132834 217242 133348
rect 248952 133320 252374 133376
rect 252430 133320 252435 133376
rect 248952 133318 252435 133320
rect 252369 133315 252435 133318
rect 307661 133242 307727 133245
rect 324313 133242 324379 133245
rect 307661 133240 310040 133242
rect 307661 133184 307666 133240
rect 307722 133184 310040 133240
rect 307661 133182 310040 133184
rect 321908 133240 324379 133242
rect 321908 133184 324318 133240
rect 324374 133184 324379 133240
rect 321908 133182 324379 133184
rect 307661 133179 307727 133182
rect 324313 133179 324379 133182
rect 252185 132834 252251 132837
rect 214005 132832 217242 132834
rect 214005 132776 214010 132832
rect 214066 132776 217242 132832
rect 214005 132774 217242 132776
rect 248952 132832 252251 132834
rect 248952 132776 252190 132832
rect 252246 132776 252251 132832
rect 248952 132774 252251 132776
rect 214005 132771 214071 132774
rect 252185 132771 252251 132774
rect 307201 132698 307267 132701
rect 307201 132696 310040 132698
rect 213913 132562 213979 132565
rect 213913 132560 216874 132562
rect 213913 132504 213918 132560
rect 213974 132510 216874 132560
rect 217366 132510 217426 132668
rect 307201 132640 307206 132696
rect 307262 132640 310040 132696
rect 307201 132638 310040 132640
rect 307201 132635 307267 132638
rect 213974 132504 217426 132510
rect 213913 132502 217426 132504
rect 213913 132499 213979 132502
rect 216814 132450 217426 132502
rect 252369 132426 252435 132429
rect 324313 132426 324379 132429
rect 248952 132424 252435 132426
rect 248952 132368 252374 132424
rect 252430 132368 252435 132424
rect 248952 132366 252435 132368
rect 321908 132424 324379 132426
rect 321908 132368 324318 132424
rect 324374 132368 324379 132424
rect 321908 132366 324379 132368
rect 252369 132363 252435 132366
rect 324313 132363 324379 132366
rect 307385 132290 307451 132293
rect 307385 132288 310040 132290
rect 307385 132232 307390 132288
rect 307446 132232 310040 132288
rect 307385 132230 310040 132232
rect 307385 132227 307451 132230
rect 214005 131474 214071 131477
rect 217182 131474 217242 131988
rect 252461 131882 252527 131885
rect 248952 131880 252527 131882
rect 248952 131824 252466 131880
rect 252522 131824 252527 131880
rect 248952 131822 252527 131824
rect 252461 131819 252527 131822
rect 307569 131882 307635 131885
rect 307569 131880 310040 131882
rect 307569 131824 307574 131880
rect 307630 131824 310040 131880
rect 307569 131822 310040 131824
rect 307569 131819 307635 131822
rect 324405 131746 324471 131749
rect 321908 131744 324471 131746
rect 321908 131688 324410 131744
rect 324466 131688 324471 131744
rect 321908 131686 324471 131688
rect 324405 131683 324471 131686
rect 252277 131474 252343 131477
rect 214005 131472 217242 131474
rect 214005 131416 214010 131472
rect 214066 131416 217242 131472
rect 214005 131414 217242 131416
rect 248952 131472 252343 131474
rect 248952 131416 252282 131472
rect 252338 131416 252343 131472
rect 248952 131414 252343 131416
rect 214005 131411 214071 131414
rect 252277 131411 252343 131414
rect 307661 131474 307727 131477
rect 307661 131472 310040 131474
rect 307661 131416 307666 131472
rect 307722 131416 310040 131472
rect 307661 131414 310040 131416
rect 307661 131411 307727 131414
rect 213913 131202 213979 131205
rect 213913 131200 216874 131202
rect 213913 131144 213918 131200
rect 213974 131144 216874 131200
rect 213913 131142 216874 131144
rect 213913 131139 213979 131142
rect 216814 131066 216874 131142
rect 217366 131066 217426 131308
rect 216814 131006 217426 131066
rect 307661 131066 307727 131069
rect 307661 131064 310040 131066
rect 307661 131008 307666 131064
rect 307722 131008 310040 131064
rect 307661 131006 310040 131008
rect 307661 131003 307727 131006
rect 251950 130930 251956 130932
rect 248952 130870 251956 130930
rect 251950 130868 251956 130870
rect 252020 130868 252026 130932
rect 324313 130930 324379 130933
rect 321908 130928 324379 130930
rect 321908 130872 324318 130928
rect 324374 130872 324379 130928
rect 321908 130870 324379 130872
rect 324313 130867 324379 130870
rect 214005 130114 214071 130117
rect 217182 130114 217242 130628
rect 309550 130554 310132 130614
rect 252461 130522 252527 130525
rect 248952 130520 252527 130522
rect 248952 130464 252466 130520
rect 252522 130464 252527 130520
rect 248952 130462 252527 130464
rect 252461 130459 252527 130462
rect 252277 130114 252343 130117
rect 214005 130112 217242 130114
rect 214005 130056 214010 130112
rect 214066 130056 217242 130112
rect 214005 130054 217242 130056
rect 248952 130112 252343 130114
rect 248952 130056 252282 130112
rect 252338 130056 252343 130112
rect 248952 130054 252343 130056
rect 214005 130051 214071 130054
rect 252277 130051 252343 130054
rect 305494 130052 305500 130116
rect 305564 130114 305570 130116
rect 309550 130114 309610 130554
rect 305564 130054 309610 130114
rect 309734 130146 310132 130206
rect 305564 130052 305570 130054
rect 307569 129978 307635 129981
rect 309734 129978 309794 130146
rect 324405 130114 324471 130117
rect 321908 130112 324471 130114
rect 321908 130056 324410 130112
rect 324466 130056 324471 130112
rect 321908 130054 324471 130056
rect 324405 130051 324471 130054
rect 307569 129976 309794 129978
rect 213913 129842 213979 129845
rect 213913 129840 216874 129842
rect 213913 129784 213918 129840
rect 213974 129784 216874 129840
rect 213913 129782 216874 129784
rect 213913 129779 213979 129782
rect 216814 129706 216874 129782
rect 217366 129706 217426 129948
rect 307569 129920 307574 129976
rect 307630 129920 309794 129976
rect 307569 129918 309794 129920
rect 307569 129915 307635 129918
rect 307477 129842 307543 129845
rect 307477 129840 310040 129842
rect 307477 129784 307482 129840
rect 307538 129784 310040 129840
rect 307477 129782 310040 129784
rect 307477 129779 307543 129782
rect 216814 129646 217426 129706
rect 252369 129570 252435 129573
rect 248952 129568 252435 129570
rect 248952 129512 252374 129568
rect 252430 129512 252435 129568
rect 248952 129510 252435 129512
rect 252369 129507 252435 129510
rect 324313 129434 324379 129437
rect 321908 129432 324379 129434
rect 321908 129376 324318 129432
rect 324374 129376 324379 129432
rect 321908 129374 324379 129376
rect 324313 129371 324379 129374
rect 66161 129298 66227 129301
rect 68142 129298 68816 129304
rect 66161 129296 68816 129298
rect 66161 129240 66166 129296
rect 66222 129244 68816 129296
rect 307569 129298 307635 129301
rect 307569 129296 310040 129298
rect 66222 129240 68202 129244
rect 66161 129238 68202 129240
rect 66161 129235 66227 129238
rect 213913 128890 213979 128893
rect 217182 128890 217242 129268
rect 307569 129240 307574 129296
rect 307630 129240 310040 129296
rect 307569 129238 310040 129240
rect 307569 129235 307635 129238
rect 252461 129162 252527 129165
rect 248952 129160 252527 129162
rect 248952 129104 252466 129160
rect 252522 129104 252527 129160
rect 248952 129102 252527 129104
rect 252461 129099 252527 129102
rect 213913 128888 217242 128890
rect 213913 128832 213918 128888
rect 213974 128832 217242 128888
rect 213913 128830 217242 128832
rect 306741 128890 306807 128893
rect 306741 128888 310040 128890
rect 306741 128832 306746 128888
rect 306802 128832 310040 128888
rect 306741 128830 310040 128832
rect 213913 128827 213979 128830
rect 306741 128827 306807 128830
rect 170254 128556 170260 128620
rect 170324 128618 170330 128620
rect 170324 128558 200130 128618
rect 170324 128556 170330 128558
rect 200070 128482 200130 128558
rect 217366 128482 217426 128724
rect 252277 128618 252343 128621
rect 324405 128618 324471 128621
rect 248952 128616 252343 128618
rect 248952 128560 252282 128616
rect 252338 128560 252343 128616
rect 248952 128558 252343 128560
rect 321908 128616 324471 128618
rect 321908 128560 324410 128616
rect 324466 128560 324471 128616
rect 321908 128558 324471 128560
rect 252277 128555 252343 128558
rect 324405 128555 324471 128558
rect 200070 128422 217426 128482
rect 307661 128482 307727 128485
rect 307661 128480 310040 128482
rect 307661 128424 307666 128480
rect 307722 128424 310040 128480
rect 307661 128422 310040 128424
rect 307661 128419 307727 128422
rect 252461 128210 252527 128213
rect 248952 128208 252527 128210
rect 248952 128152 252466 128208
rect 252522 128152 252527 128208
rect 248952 128150 252527 128152
rect 252461 128147 252527 128150
rect 67541 128074 67607 128077
rect 68142 128074 68816 128080
rect 67541 128072 68816 128074
rect 67541 128016 67546 128072
rect 67602 128020 68816 128072
rect 307477 128074 307543 128077
rect 307477 128072 310040 128074
rect 67602 128016 68202 128020
rect 67541 128014 68202 128016
rect 67541 128011 67607 128014
rect 213453 127530 213519 127533
rect 217182 127530 217242 128044
rect 307477 128016 307482 128072
rect 307538 128016 310040 128072
rect 307477 128014 310040 128016
rect 307477 128011 307543 128014
rect 324313 127802 324379 127805
rect 321908 127800 324379 127802
rect 321908 127744 324318 127800
rect 324374 127744 324379 127800
rect 321908 127742 324379 127744
rect 324313 127739 324379 127742
rect 252369 127666 252435 127669
rect 248952 127664 252435 127666
rect 248952 127608 252374 127664
rect 252430 127608 252435 127664
rect 248952 127606 252435 127608
rect 252369 127603 252435 127606
rect 307569 127666 307635 127669
rect 307569 127664 310040 127666
rect 307569 127608 307574 127664
rect 307630 127608 310040 127664
rect 307569 127606 310040 127608
rect 307569 127603 307635 127606
rect 213453 127528 217242 127530
rect 213453 127472 213458 127528
rect 213514 127472 217242 127528
rect 213453 127470 217242 127472
rect 321645 127530 321711 127533
rect 321645 127528 321754 127530
rect 321645 127472 321650 127528
rect 321706 127472 321754 127528
rect 213453 127467 213519 127470
rect 321645 127467 321754 127472
rect 173014 127196 173020 127260
rect 173084 127258 173090 127260
rect 173084 127198 213746 127258
rect 173084 127196 173090 127198
rect 169150 127060 169156 127124
rect 169220 127122 169226 127124
rect 213453 127122 213519 127125
rect 169220 127120 213519 127122
rect 169220 127064 213458 127120
rect 213514 127064 213519 127120
rect 169220 127062 213519 127064
rect 213686 127122 213746 127198
rect 217366 127122 217426 127364
rect 252461 127258 252527 127261
rect 248952 127256 252527 127258
rect 248952 127200 252466 127256
rect 252522 127200 252527 127256
rect 248952 127198 252527 127200
rect 252461 127195 252527 127198
rect 307661 127258 307727 127261
rect 307661 127256 310040 127258
rect 307661 127200 307666 127256
rect 307722 127200 310040 127256
rect 307661 127198 310040 127200
rect 307661 127195 307727 127198
rect 213686 127062 217426 127122
rect 321694 127092 321754 127467
rect 169220 127060 169226 127062
rect 213453 127059 213519 127062
rect 307477 126850 307543 126853
rect 307477 126848 310040 126850
rect 307477 126792 307482 126848
rect 307538 126792 310040 126848
rect 307477 126790 310040 126792
rect 307477 126787 307543 126790
rect 252461 126714 252527 126717
rect 248952 126712 252527 126714
rect 65149 126306 65215 126309
rect 68142 126306 68816 126312
rect 65149 126304 68816 126306
rect 65149 126248 65154 126304
rect 65210 126252 68816 126304
rect 65210 126248 68202 126252
rect 65149 126246 68202 126248
rect 65149 126243 65215 126246
rect 214005 126170 214071 126173
rect 217182 126170 217242 126684
rect 248952 126656 252466 126712
rect 252522 126656 252527 126712
rect 248952 126654 252527 126656
rect 252461 126651 252527 126654
rect 307569 126442 307635 126445
rect 307569 126440 310040 126442
rect 307569 126384 307574 126440
rect 307630 126384 310040 126440
rect 307569 126382 310040 126384
rect 307569 126379 307635 126382
rect 251909 126306 251975 126309
rect 324313 126306 324379 126309
rect 248952 126304 251975 126306
rect 248952 126248 251914 126304
rect 251970 126248 251975 126304
rect 248952 126246 251975 126248
rect 321908 126304 324379 126306
rect 321908 126248 324318 126304
rect 324374 126248 324379 126304
rect 321908 126246 324379 126248
rect 251909 126243 251975 126246
rect 324313 126243 324379 126246
rect 214005 126168 217242 126170
rect 214005 126112 214010 126168
rect 214066 126112 217242 126168
rect 214005 126110 217242 126112
rect 214005 126107 214071 126110
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 213913 125762 213979 125765
rect 217182 125762 217242 126004
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 307661 125898 307727 125901
rect 307661 125896 310040 125898
rect 307661 125840 307666 125896
rect 307722 125840 310040 125896
rect 583520 125884 584960 125974
rect 307661 125838 310040 125840
rect 307661 125835 307727 125838
rect 252369 125762 252435 125765
rect 213913 125760 217242 125762
rect 213913 125704 213918 125760
rect 213974 125704 217242 125760
rect 213913 125702 217242 125704
rect 248952 125760 252435 125762
rect 248952 125704 252374 125760
rect 252430 125704 252435 125760
rect 248952 125702 252435 125704
rect 213913 125699 213979 125702
rect 252369 125699 252435 125702
rect 307569 125490 307635 125493
rect 324957 125490 325023 125493
rect 307569 125488 310040 125490
rect 307569 125432 307574 125488
rect 307630 125432 310040 125488
rect 307569 125430 310040 125432
rect 321908 125488 325023 125490
rect 321908 125432 324962 125488
rect 325018 125432 325023 125488
rect 321908 125430 325023 125432
rect 307569 125427 307635 125430
rect 324957 125427 325023 125430
rect 252369 125354 252435 125357
rect 248952 125352 252435 125354
rect 66069 125218 66135 125221
rect 68142 125218 68816 125224
rect 66069 125216 68816 125218
rect 66069 125160 66074 125216
rect 66130 125164 68816 125216
rect 66130 125160 68202 125164
rect 66069 125158 68202 125160
rect 66069 125155 66135 125158
rect 214005 124810 214071 124813
rect 217182 124810 217242 125324
rect 248952 125296 252374 125352
rect 252430 125296 252435 125352
rect 248952 125294 252435 125296
rect 252369 125291 252435 125294
rect 306925 125082 306991 125085
rect 306925 125080 310040 125082
rect 306925 125024 306930 125080
rect 306986 125024 310040 125080
rect 306925 125022 310040 125024
rect 306925 125019 306991 125022
rect 252461 124810 252527 124813
rect 325601 124810 325667 124813
rect 214005 124808 217242 124810
rect 214005 124752 214010 124808
rect 214066 124752 217242 124808
rect 214005 124750 217242 124752
rect 248952 124808 252527 124810
rect 248952 124752 252466 124808
rect 252522 124752 252527 124808
rect 248952 124750 252527 124752
rect 321908 124808 325667 124810
rect 321908 124752 325606 124808
rect 325662 124752 325667 124808
rect 321908 124750 325667 124752
rect 214005 124747 214071 124750
rect 252461 124747 252527 124750
rect 325601 124747 325667 124750
rect 307293 124674 307359 124677
rect 307293 124672 310040 124674
rect 213913 124402 213979 124405
rect 217182 124402 217242 124644
rect 307293 124616 307298 124672
rect 307354 124616 310040 124672
rect 307293 124614 310040 124616
rect 307293 124611 307359 124614
rect 252185 124402 252251 124405
rect 213913 124400 217242 124402
rect 213913 124344 213918 124400
rect 213974 124344 217242 124400
rect 213913 124342 217242 124344
rect 248952 124400 252251 124402
rect 248952 124344 252190 124400
rect 252246 124344 252251 124400
rect 248952 124342 252251 124344
rect 213913 124339 213979 124342
rect 252185 124339 252251 124342
rect 307661 124266 307727 124269
rect 321553 124266 321619 124269
rect 307661 124264 310040 124266
rect 307661 124208 307666 124264
rect 307722 124208 310040 124264
rect 307661 124206 310040 124208
rect 321510 124264 321619 124266
rect 321510 124208 321558 124264
rect 321614 124208 321619 124264
rect 307661 124203 307727 124206
rect 321510 124203 321619 124208
rect -960 123572 480 123812
rect 65977 123586 66043 123589
rect 68142 123586 68816 123592
rect 65977 123584 68816 123586
rect 65977 123528 65982 123584
rect 66038 123532 68816 123584
rect 213913 123586 213979 123589
rect 217182 123586 217242 124100
rect 252277 123994 252343 123997
rect 248952 123992 252343 123994
rect 248952 123936 252282 123992
rect 252338 123936 252343 123992
rect 321510 123964 321570 124203
rect 248952 123934 252343 123936
rect 252277 123931 252343 123934
rect 307477 123858 307543 123861
rect 307477 123856 310040 123858
rect 307477 123800 307482 123856
rect 307538 123800 310040 123856
rect 307477 123798 310040 123800
rect 307477 123795 307543 123798
rect 213913 123584 217242 123586
rect 66038 123528 68202 123532
rect 65977 123526 68202 123528
rect 213913 123528 213918 123584
rect 213974 123528 217242 123584
rect 213913 123526 217242 123528
rect 65977 123523 66043 123526
rect 213913 123523 213979 123526
rect 252461 123450 252527 123453
rect 248952 123448 252527 123450
rect 64781 122906 64847 122909
rect 65977 122906 66043 122909
rect 64781 122904 66043 122906
rect 64781 122848 64786 122904
rect 64842 122848 65982 122904
rect 66038 122848 66043 122904
rect 64781 122846 66043 122848
rect 64781 122843 64847 122846
rect 65977 122843 66043 122846
rect 213913 122906 213979 122909
rect 217182 122906 217242 123420
rect 248952 123392 252466 123448
rect 252522 123392 252527 123448
rect 248952 123390 252527 123392
rect 252461 123387 252527 123390
rect 307661 123450 307727 123453
rect 307661 123448 310040 123450
rect 307661 123392 307666 123448
rect 307722 123392 310040 123448
rect 307661 123390 310040 123392
rect 307661 123387 307727 123390
rect 324313 123178 324379 123181
rect 321908 123176 324379 123178
rect 321908 123120 324318 123176
rect 324374 123120 324379 123176
rect 321908 123118 324379 123120
rect 324313 123115 324379 123118
rect 252369 123042 252435 123045
rect 248952 123040 252435 123042
rect 248952 122984 252374 123040
rect 252430 122984 252435 123040
rect 248952 122982 252435 122984
rect 252369 122979 252435 122982
rect 307569 123042 307635 123045
rect 307569 123040 310040 123042
rect 307569 122984 307574 123040
rect 307630 122984 310040 123040
rect 307569 122982 310040 122984
rect 307569 122979 307635 122982
rect 213913 122904 217242 122906
rect 213913 122848 213918 122904
rect 213974 122848 217242 122904
rect 213913 122846 217242 122848
rect 213913 122843 213979 122846
rect 65977 122634 66043 122637
rect 68142 122634 68816 122640
rect 65977 122632 68816 122634
rect 65977 122576 65982 122632
rect 66038 122580 68816 122632
rect 66038 122576 68202 122580
rect 65977 122574 68202 122576
rect 65977 122571 66043 122574
rect 214005 122226 214071 122229
rect 217182 122226 217242 122740
rect 252461 122498 252527 122501
rect 248952 122496 252527 122498
rect 248952 122440 252466 122496
rect 252522 122440 252527 122496
rect 248952 122438 252527 122440
rect 252461 122435 252527 122438
rect 307477 122498 307543 122501
rect 324313 122498 324379 122501
rect 307477 122496 310040 122498
rect 307477 122440 307482 122496
rect 307538 122440 310040 122496
rect 307477 122438 310040 122440
rect 321908 122496 324379 122498
rect 321908 122440 324318 122496
rect 324374 122440 324379 122496
rect 321908 122438 324379 122440
rect 307477 122435 307543 122438
rect 324313 122435 324379 122438
rect 214005 122224 217242 122226
rect 214005 122168 214010 122224
rect 214066 122168 217242 122224
rect 214005 122166 217242 122168
rect 214005 122163 214071 122166
rect 253197 122090 253263 122093
rect 248952 122088 253263 122090
rect 213913 121818 213979 121821
rect 217182 121818 217242 122060
rect 248952 122032 253202 122088
rect 253258 122032 253263 122088
rect 248952 122030 253263 122032
rect 253197 122027 253263 122030
rect 307569 122090 307635 122093
rect 307569 122088 310040 122090
rect 307569 122032 307574 122088
rect 307630 122032 310040 122088
rect 307569 122030 310040 122032
rect 307569 122027 307635 122030
rect 213913 121816 217242 121818
rect 213913 121760 213918 121816
rect 213974 121760 217242 121816
rect 213913 121758 217242 121760
rect 213913 121755 213979 121758
rect 307661 121682 307727 121685
rect 323117 121682 323183 121685
rect 307661 121680 310040 121682
rect 307661 121624 307666 121680
rect 307722 121624 310040 121680
rect 307661 121622 310040 121624
rect 321908 121680 323183 121682
rect 321908 121624 323122 121680
rect 323178 121624 323183 121680
rect 321908 121622 323183 121624
rect 307661 121619 307727 121622
rect 323117 121619 323183 121622
rect 252369 121546 252435 121549
rect 248952 121544 252435 121546
rect 248952 121488 252374 121544
rect 252430 121488 252435 121544
rect 248952 121486 252435 121488
rect 252369 121483 252435 121486
rect 67449 120866 67515 120869
rect 68142 120866 68816 120872
rect 67449 120864 68816 120866
rect 67449 120808 67454 120864
rect 67510 120812 68816 120864
rect 213913 120866 213979 120869
rect 217182 120866 217242 121380
rect 307477 121274 307543 121277
rect 307477 121272 310040 121274
rect 307477 121216 307482 121272
rect 307538 121216 310040 121272
rect 307477 121214 310040 121216
rect 307477 121211 307543 121214
rect 252461 121138 252527 121141
rect 248952 121136 252527 121138
rect 248952 121080 252466 121136
rect 252522 121080 252527 121136
rect 248952 121078 252527 121080
rect 252461 121075 252527 121078
rect 213913 120864 217242 120866
rect 67510 120808 68202 120812
rect 67449 120806 68202 120808
rect 213913 120808 213918 120864
rect 213974 120808 217242 120864
rect 213913 120806 217242 120808
rect 307569 120866 307635 120869
rect 324313 120866 324379 120869
rect 307569 120864 310040 120866
rect 307569 120808 307574 120864
rect 307630 120808 310040 120864
rect 307569 120806 310040 120808
rect 321908 120864 324379 120866
rect 321908 120808 324318 120864
rect 324374 120808 324379 120864
rect 321908 120806 324379 120808
rect 67449 120803 67515 120806
rect 213913 120803 213979 120806
rect 307569 120803 307635 120806
rect 324313 120803 324379 120806
rect 213269 120186 213335 120189
rect 217182 120186 217242 120700
rect 252369 120594 252435 120597
rect 248952 120592 252435 120594
rect 248952 120536 252374 120592
rect 252430 120536 252435 120592
rect 248952 120534 252435 120536
rect 252369 120531 252435 120534
rect 307661 120458 307727 120461
rect 307661 120456 310040 120458
rect 307661 120400 307666 120456
rect 307722 120400 310040 120456
rect 307661 120398 310040 120400
rect 307661 120395 307727 120398
rect 252277 120186 252343 120189
rect 324405 120186 324471 120189
rect 213269 120184 217242 120186
rect 213269 120128 213274 120184
rect 213330 120128 217242 120184
rect 213269 120126 217242 120128
rect 248952 120184 252343 120186
rect 248952 120128 252282 120184
rect 252338 120128 252343 120184
rect 248952 120126 252343 120128
rect 321908 120184 324471 120186
rect 321908 120128 324410 120184
rect 324466 120128 324471 120184
rect 321908 120126 324471 120128
rect 213269 120123 213335 120126
rect 252277 120123 252343 120126
rect 324405 120123 324471 120126
rect 307477 120050 307543 120053
rect 307477 120048 310040 120050
rect 214005 119642 214071 119645
rect 217182 119642 217242 120020
rect 307477 119992 307482 120048
rect 307538 119992 310040 120048
rect 307477 119990 310040 119992
rect 307477 119987 307543 119990
rect 252461 119642 252527 119645
rect 214005 119640 217242 119642
rect 214005 119584 214010 119640
rect 214066 119584 217242 119640
rect 214005 119582 217242 119584
rect 248952 119640 252527 119642
rect 248952 119584 252466 119640
rect 252522 119584 252527 119640
rect 248952 119582 252527 119584
rect 214005 119579 214071 119582
rect 252461 119579 252527 119582
rect 307569 119642 307635 119645
rect 307569 119640 310040 119642
rect 307569 119584 307574 119640
rect 307630 119584 310040 119640
rect 307569 119582 310040 119584
rect 307569 119579 307635 119582
rect 214097 119098 214163 119101
rect 217182 119098 217242 119476
rect 324313 119370 324379 119373
rect 321908 119368 324379 119370
rect 321908 119312 324318 119368
rect 324374 119312 324379 119368
rect 321908 119310 324379 119312
rect 324313 119307 324379 119310
rect 252461 119234 252527 119237
rect 248952 119232 252527 119234
rect 248952 119176 252466 119232
rect 252522 119176 252527 119232
rect 248952 119174 252527 119176
rect 252461 119171 252527 119174
rect 214097 119096 217242 119098
rect 214097 119040 214102 119096
rect 214158 119040 217242 119096
rect 214097 119038 217242 119040
rect 307661 119098 307727 119101
rect 307661 119096 310040 119098
rect 307661 119040 307666 119096
rect 307722 119040 310040 119096
rect 307661 119038 310040 119040
rect 214097 119035 214163 119038
rect 307661 119035 307727 119038
rect 213913 118962 213979 118965
rect 213913 118960 217242 118962
rect 213913 118904 213918 118960
rect 213974 118904 217242 118960
rect 213913 118902 217242 118904
rect 213913 118899 213979 118902
rect 217182 118796 217242 118902
rect 252369 118826 252435 118829
rect 248952 118824 252435 118826
rect 248952 118768 252374 118824
rect 252430 118768 252435 118824
rect 248952 118766 252435 118768
rect 252369 118763 252435 118766
rect 305821 118826 305887 118829
rect 307569 118826 307635 118829
rect 305821 118824 307635 118826
rect 305821 118768 305826 118824
rect 305882 118768 307574 118824
rect 307630 118768 307635 118824
rect 305821 118766 307635 118768
rect 305821 118763 305887 118766
rect 307569 118763 307635 118766
rect 306557 118690 306623 118693
rect 306557 118688 310040 118690
rect 306557 118632 306562 118688
rect 306618 118632 310040 118688
rect 306557 118630 310040 118632
rect 306557 118627 306623 118630
rect 324313 118554 324379 118557
rect 321908 118552 324379 118554
rect 321908 118496 324318 118552
rect 324374 118496 324379 118552
rect 321908 118494 324379 118496
rect 324313 118491 324379 118494
rect 252461 118282 252527 118285
rect 248952 118280 252527 118282
rect 248952 118224 252466 118280
rect 252522 118224 252527 118280
rect 248952 118222 252527 118224
rect 252461 118219 252527 118222
rect 309550 118178 310132 118238
rect 213361 117602 213427 117605
rect 217182 117602 217242 118116
rect 299974 118084 299980 118148
rect 300044 118146 300050 118148
rect 309550 118146 309610 118178
rect 300044 118086 309610 118146
rect 300044 118084 300050 118086
rect 252369 117874 252435 117877
rect 248952 117872 252435 117874
rect 248952 117816 252374 117872
rect 252430 117816 252435 117872
rect 248952 117814 252435 117816
rect 252369 117811 252435 117814
rect 307569 117874 307635 117877
rect 324405 117874 324471 117877
rect 307569 117872 310040 117874
rect 307569 117816 307574 117872
rect 307630 117816 310040 117872
rect 307569 117814 310040 117816
rect 321908 117872 324471 117874
rect 321908 117816 324410 117872
rect 324466 117816 324471 117872
rect 321908 117814 324471 117816
rect 307569 117811 307635 117814
rect 324405 117811 324471 117814
rect 213361 117600 217242 117602
rect 213361 117544 213366 117600
rect 213422 117544 217242 117600
rect 213361 117542 217242 117544
rect 213361 117539 213427 117542
rect 307661 117466 307727 117469
rect 307661 117464 310040 117466
rect 213913 117330 213979 117333
rect 213913 117328 216874 117330
rect 213913 117272 213918 117328
rect 213974 117272 216874 117328
rect 213913 117270 216874 117272
rect 213913 117267 213979 117270
rect 216814 117194 216874 117270
rect 217366 117194 217426 117436
rect 307661 117408 307666 117464
rect 307722 117408 310040 117464
rect 307661 117406 310040 117408
rect 307661 117403 307727 117406
rect 251633 117330 251699 117333
rect 248952 117328 251699 117330
rect 248952 117272 251638 117328
rect 251694 117272 251699 117328
rect 248952 117270 251699 117272
rect 251633 117267 251699 117270
rect 216814 117134 217426 117194
rect 307569 117058 307635 117061
rect 307569 117056 310040 117058
rect 307569 117000 307574 117056
rect 307630 117000 310040 117056
rect 307569 116998 310040 117000
rect 307569 116995 307635 116998
rect 252001 116922 252067 116925
rect 248952 116920 252067 116922
rect 248952 116864 252006 116920
rect 252062 116864 252067 116920
rect 248952 116862 252067 116864
rect 252001 116859 252067 116862
rect 214005 116242 214071 116245
rect 217182 116242 217242 116756
rect 306741 116650 306807 116653
rect 306741 116648 310040 116650
rect 306741 116592 306746 116648
rect 306802 116592 310040 116648
rect 306741 116590 310040 116592
rect 306741 116587 306807 116590
rect 321878 116514 321938 117028
rect 321878 116454 325710 116514
rect 252461 116378 252527 116381
rect 324313 116378 324379 116381
rect 248952 116376 252527 116378
rect 248952 116320 252466 116376
rect 252522 116320 252527 116376
rect 248952 116318 252527 116320
rect 321908 116376 324379 116378
rect 321908 116320 324318 116376
rect 324374 116320 324379 116376
rect 321908 116318 324379 116320
rect 252461 116315 252527 116318
rect 324313 116315 324379 116318
rect 214005 116240 217242 116242
rect 214005 116184 214010 116240
rect 214066 116184 217242 116240
rect 214005 116182 217242 116184
rect 307661 116242 307727 116245
rect 307661 116240 310040 116242
rect 307661 116184 307666 116240
rect 307722 116184 310040 116240
rect 307661 116182 310040 116184
rect 214005 116179 214071 116182
rect 307661 116179 307727 116182
rect 213913 115970 213979 115973
rect 213913 115968 216874 115970
rect 213913 115912 213918 115968
rect 213974 115912 216874 115968
rect 213913 115910 216874 115912
rect 213913 115907 213979 115910
rect 166901 115836 166967 115837
rect 166901 115834 166948 115836
rect 166856 115832 166948 115834
rect 166856 115776 166906 115832
rect 166856 115774 166948 115776
rect 166901 115772 166948 115774
rect 167012 115772 167018 115836
rect 216814 115834 216874 115910
rect 217366 115834 217426 116076
rect 252461 115970 252527 115973
rect 248952 115968 252527 115970
rect 248952 115912 252466 115968
rect 252522 115912 252527 115968
rect 248952 115910 252527 115912
rect 325650 115970 325710 116454
rect 335486 115970 335492 115972
rect 325650 115910 335492 115970
rect 252461 115907 252527 115910
rect 335486 115908 335492 115910
rect 335556 115908 335562 115972
rect 216814 115774 217426 115834
rect 166901 115771 166967 115772
rect 307477 115698 307543 115701
rect 307477 115696 310040 115698
rect 307477 115640 307482 115696
rect 307538 115640 310040 115696
rect 307477 115638 310040 115640
rect 307477 115635 307543 115638
rect 252277 115426 252343 115429
rect 248952 115424 252343 115426
rect 214005 115018 214071 115021
rect 217182 115018 217242 115396
rect 248952 115368 252282 115424
rect 252338 115368 252343 115424
rect 248952 115366 252343 115368
rect 252277 115363 252343 115366
rect 307569 115290 307635 115293
rect 307569 115288 310040 115290
rect 307569 115232 307574 115288
rect 307630 115232 310040 115288
rect 307569 115230 310040 115232
rect 307569 115227 307635 115230
rect 252369 115018 252435 115021
rect 214005 115016 217242 115018
rect 214005 114960 214010 115016
rect 214066 114960 217242 115016
rect 214005 114958 217242 114960
rect 248952 115016 252435 115018
rect 248952 114960 252374 115016
rect 252430 114960 252435 115016
rect 248952 114958 252435 114960
rect 321878 115018 321938 115532
rect 323485 115018 323551 115021
rect 321878 115016 323551 115018
rect 321878 114960 323490 115016
rect 323546 114960 323551 115016
rect 321878 114958 323551 114960
rect 214005 114955 214071 114958
rect 252369 114955 252435 114958
rect 323485 114955 323551 114958
rect 307661 114882 307727 114885
rect 307661 114880 310040 114882
rect 213913 114610 213979 114613
rect 217366 114610 217426 114852
rect 307661 114824 307666 114880
rect 307722 114824 310040 114880
rect 307661 114822 310040 114824
rect 307661 114819 307727 114822
rect 331438 114746 331444 114748
rect 321908 114686 331444 114746
rect 331438 114684 331444 114686
rect 331508 114684 331514 114748
rect 213913 114608 217426 114610
rect 213913 114552 213918 114608
rect 213974 114552 217426 114608
rect 213913 114550 217426 114552
rect 323485 114610 323551 114613
rect 345054 114610 345060 114612
rect 323485 114608 345060 114610
rect 323485 114552 323490 114608
rect 323546 114552 345060 114608
rect 323485 114550 345060 114552
rect 213913 114547 213979 114550
rect 323485 114547 323551 114550
rect 345054 114548 345060 114550
rect 345124 114548 345130 114612
rect 252461 114474 252527 114477
rect 248952 114472 252527 114474
rect 248952 114416 252466 114472
rect 252522 114416 252527 114472
rect 248952 114414 252527 114416
rect 252461 114411 252527 114414
rect 309133 114474 309199 114477
rect 309133 114472 310040 114474
rect 309133 114416 309138 114472
rect 309194 114416 310040 114472
rect 309133 114414 310040 114416
rect 309133 114411 309199 114414
rect 213913 113658 213979 113661
rect 217182 113658 217242 114172
rect 252369 114066 252435 114069
rect 248952 114064 252435 114066
rect 248952 114008 252374 114064
rect 252430 114008 252435 114064
rect 248952 114006 252435 114008
rect 252369 114003 252435 114006
rect 307150 114004 307156 114068
rect 307220 114066 307226 114068
rect 324313 114066 324379 114069
rect 307220 114006 310040 114066
rect 321908 114064 324379 114066
rect 321908 114008 324318 114064
rect 324374 114008 324379 114064
rect 321908 114006 324379 114008
rect 307220 114004 307226 114006
rect 324313 114003 324379 114006
rect 213913 113656 217242 113658
rect 213913 113600 213918 113656
rect 213974 113600 217242 113656
rect 213913 113598 217242 113600
rect 307661 113658 307727 113661
rect 307661 113656 310040 113658
rect 307661 113600 307666 113656
rect 307722 113600 310040 113656
rect 307661 113598 310040 113600
rect 213913 113595 213979 113598
rect 307661 113595 307727 113598
rect 252277 113522 252343 113525
rect 248952 113520 252343 113522
rect 214005 113250 214071 113253
rect 217366 113250 217426 113492
rect 248952 113464 252282 113520
rect 252338 113464 252343 113520
rect 248952 113462 252343 113464
rect 252277 113459 252343 113462
rect 301814 113460 301820 113524
rect 301884 113522 301890 113524
rect 301884 113462 309380 113522
rect 301884 113460 301890 113462
rect 214005 113248 217426 113250
rect 214005 113192 214010 113248
rect 214066 113192 217426 113248
rect 214005 113190 217426 113192
rect 307569 113250 307635 113253
rect 309320 113250 309380 113462
rect 324405 113250 324471 113253
rect 307569 113248 309150 113250
rect 307569 113192 307574 113248
rect 307630 113192 309150 113248
rect 307569 113190 309150 113192
rect 309320 113190 310040 113250
rect 321908 113248 324471 113250
rect 321908 113192 324410 113248
rect 324466 113192 324471 113248
rect 321908 113190 324471 113192
rect 214005 113187 214071 113190
rect 307569 113187 307635 113190
rect 309090 113117 309150 113190
rect 324405 113187 324471 113190
rect 309090 113112 309199 113117
rect 248860 113010 249442 113070
rect 309090 113056 309138 113112
rect 309194 113056 309199 113112
rect 309090 113054 309199 113056
rect 309133 113051 309199 113054
rect 249382 112978 249442 113010
rect 258574 112978 258580 112980
rect 249382 112918 258580 112978
rect 258574 112916 258580 112918
rect 258644 112916 258650 112980
rect 582741 112842 582807 112845
rect 583520 112842 584960 112932
rect 582741 112840 584960 112842
rect 214005 112298 214071 112301
rect 217182 112298 217242 112812
rect 582741 112784 582746 112840
rect 582802 112784 584960 112840
rect 582741 112782 584960 112784
rect 582741 112779 582807 112782
rect 251766 112706 251772 112708
rect 248952 112646 251772 112706
rect 251766 112644 251772 112646
rect 251836 112644 251842 112708
rect 583520 112692 584960 112782
rect 214005 112296 217242 112298
rect 214005 112240 214010 112296
rect 214066 112240 217242 112296
rect 214005 112238 217242 112240
rect 309550 112602 310132 112662
rect 214005 112235 214071 112238
rect 252461 112162 252527 112165
rect 248952 112160 252527 112162
rect 213913 111890 213979 111893
rect 217182 111890 217242 112132
rect 248952 112104 252466 112160
rect 252522 112104 252527 112160
rect 248952 112102 252527 112104
rect 252461 112099 252527 112102
rect 302918 112100 302924 112164
rect 302988 112162 302994 112164
rect 309550 112162 309610 112602
rect 324313 112434 324379 112437
rect 321908 112432 324379 112434
rect 321908 112376 324318 112432
rect 324374 112376 324379 112432
rect 321908 112374 324379 112376
rect 324313 112371 324379 112374
rect 302988 112102 309610 112162
rect 309734 112194 310132 112254
rect 302988 112100 302994 112102
rect 307661 112026 307727 112029
rect 309734 112026 309794 112194
rect 307661 112024 309794 112026
rect 307661 111968 307666 112024
rect 307722 111968 309794 112024
rect 307661 111966 309794 111968
rect 307661 111963 307727 111966
rect 213913 111888 217242 111890
rect 213913 111832 213918 111888
rect 213974 111832 217242 111888
rect 213913 111830 217242 111832
rect 307477 111890 307543 111893
rect 307477 111888 310040 111890
rect 307477 111832 307482 111888
rect 307538 111832 310040 111888
rect 307477 111830 310040 111832
rect 213913 111827 213979 111830
rect 307477 111827 307543 111830
rect 168005 111754 168071 111757
rect 252369 111754 252435 111757
rect 164694 111752 168071 111754
rect 164694 111696 168010 111752
rect 168066 111696 168071 111752
rect 164694 111694 168071 111696
rect 248952 111752 252435 111754
rect 248952 111696 252374 111752
rect 252430 111696 252435 111752
rect 248952 111694 252435 111696
rect 168005 111691 168071 111694
rect 252369 111691 252435 111694
rect 307569 111482 307635 111485
rect 307569 111480 310040 111482
rect 214005 110938 214071 110941
rect 217182 110938 217242 111452
rect 307569 111424 307574 111480
rect 307630 111424 310040 111480
rect 307569 111422 310040 111424
rect 307569 111419 307635 111422
rect 252461 111210 252527 111213
rect 248952 111208 252527 111210
rect 248952 111152 252466 111208
rect 252522 111152 252527 111208
rect 248952 111150 252527 111152
rect 321878 111210 321938 111724
rect 323485 111210 323551 111213
rect 321878 111208 323551 111210
rect 321878 111152 323490 111208
rect 323546 111152 323551 111208
rect 321878 111150 323551 111152
rect 252461 111147 252527 111150
rect 323485 111147 323551 111150
rect 307661 111074 307727 111077
rect 307661 111072 310040 111074
rect 307661 111016 307666 111072
rect 307722 111016 310040 111072
rect 307661 111014 310040 111016
rect 307661 111011 307727 111014
rect 214005 110936 217242 110938
rect 214005 110880 214010 110936
rect 214066 110880 217242 110936
rect 214005 110878 217242 110880
rect 214005 110875 214071 110878
rect 251909 110802 251975 110805
rect 248952 110800 251975 110802
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 213913 110530 213979 110533
rect 217182 110530 217242 110772
rect 248952 110744 251914 110800
rect 251970 110744 251975 110800
rect 248952 110742 251975 110744
rect 251909 110739 251975 110742
rect 305637 110666 305703 110669
rect 321878 110666 321938 110908
rect 332542 110666 332548 110668
rect 305637 110664 310040 110666
rect 305637 110608 305642 110664
rect 305698 110608 310040 110664
rect 305637 110606 310040 110608
rect 321878 110606 332548 110666
rect 305637 110603 305703 110606
rect 332542 110604 332548 110606
rect 332612 110604 332618 110668
rect 213913 110528 217242 110530
rect 213913 110472 213918 110528
rect 213974 110472 217242 110528
rect 213913 110470 217242 110472
rect 323485 110530 323551 110533
rect 338246 110530 338252 110532
rect 323485 110528 338252 110530
rect 323485 110472 323490 110528
rect 323546 110472 338252 110528
rect 323485 110470 338252 110472
rect 213913 110467 213979 110470
rect 323485 110467 323551 110470
rect 338246 110468 338252 110470
rect 338316 110468 338322 110532
rect 252461 110258 252527 110261
rect 248952 110256 252527 110258
rect 168097 110122 168163 110125
rect 164694 110120 168163 110122
rect 164694 110064 168102 110120
rect 168158 110064 168163 110120
rect 164694 110062 168163 110064
rect 168097 110059 168163 110062
rect 214005 109714 214071 109717
rect 217182 109714 217242 110228
rect 248952 110200 252466 110256
rect 252522 110200 252527 110256
rect 248952 110198 252527 110200
rect 252461 110195 252527 110198
rect 307477 110258 307543 110261
rect 307477 110256 310040 110258
rect 307477 110200 307482 110256
rect 307538 110200 310040 110256
rect 307477 110198 310040 110200
rect 307477 110195 307543 110198
rect 251633 109850 251699 109853
rect 248952 109848 251699 109850
rect 248952 109792 251638 109848
rect 251694 109792 251699 109848
rect 248952 109790 251699 109792
rect 251633 109787 251699 109790
rect 307569 109850 307635 109853
rect 307569 109848 310040 109850
rect 307569 109792 307574 109848
rect 307630 109792 310040 109848
rect 307569 109790 310040 109792
rect 307569 109787 307635 109790
rect 214005 109712 217242 109714
rect 214005 109656 214010 109712
rect 214066 109656 217242 109712
rect 214005 109654 217242 109656
rect 214005 109651 214071 109654
rect 321878 109578 321938 110092
rect 334198 109578 334204 109580
rect 213913 109306 213979 109309
rect 217182 109306 217242 109548
rect 321878 109518 334204 109578
rect 334198 109516 334204 109518
rect 334268 109516 334274 109580
rect 252369 109306 252435 109309
rect 213913 109304 217242 109306
rect 213913 109248 213918 109304
rect 213974 109248 217242 109304
rect 213913 109246 217242 109248
rect 248952 109304 252435 109306
rect 248952 109248 252374 109304
rect 252430 109248 252435 109304
rect 248952 109246 252435 109248
rect 213913 109243 213979 109246
rect 252369 109243 252435 109246
rect 307661 109306 307727 109309
rect 307661 109304 310040 109306
rect 307661 109248 307666 109304
rect 307722 109248 310040 109304
rect 307661 109246 310040 109248
rect 307661 109243 307727 109246
rect 321878 109170 321938 109412
rect 335118 109170 335124 109172
rect 321878 109110 335124 109170
rect 335118 109108 335124 109110
rect 335188 109108 335194 109172
rect 252093 108898 252159 108901
rect 248952 108896 252159 108898
rect 168005 108762 168071 108765
rect 164694 108760 168071 108762
rect 164694 108704 168010 108760
rect 168066 108704 168071 108760
rect 164694 108702 168071 108704
rect 168005 108699 168071 108702
rect 214833 108354 214899 108357
rect 217182 108354 217242 108868
rect 248952 108840 252098 108896
rect 252154 108840 252159 108896
rect 248952 108838 252159 108840
rect 252093 108835 252159 108838
rect 307477 108898 307543 108901
rect 307477 108896 310040 108898
rect 307477 108840 307482 108896
rect 307538 108840 310040 108896
rect 307477 108838 310040 108840
rect 307477 108835 307543 108838
rect 324313 108626 324379 108629
rect 321908 108624 324379 108626
rect 321908 108568 324318 108624
rect 324374 108568 324379 108624
rect 321908 108566 324379 108568
rect 324313 108563 324379 108566
rect 307661 108490 307727 108493
rect 307661 108488 310040 108490
rect 307661 108432 307666 108488
rect 307722 108432 310040 108488
rect 307661 108430 310040 108432
rect 307661 108427 307727 108430
rect 252461 108354 252527 108357
rect 214833 108352 217242 108354
rect 214833 108296 214838 108352
rect 214894 108296 217242 108352
rect 214833 108294 217242 108296
rect 248952 108352 252527 108354
rect 248952 108296 252466 108352
rect 252522 108296 252527 108352
rect 248952 108294 252527 108296
rect 214833 108291 214899 108294
rect 252461 108291 252527 108294
rect 213913 107946 213979 107949
rect 217182 107946 217242 108188
rect 307569 108082 307635 108085
rect 307569 108080 310040 108082
rect 307569 108024 307574 108080
rect 307630 108024 310040 108080
rect 307569 108022 310040 108024
rect 307569 108019 307635 108022
rect 252369 107946 252435 107949
rect 213913 107944 217242 107946
rect 213913 107888 213918 107944
rect 213974 107888 217242 107944
rect 213913 107886 217242 107888
rect 248952 107944 252435 107946
rect 248952 107888 252374 107944
rect 252430 107888 252435 107944
rect 248952 107886 252435 107888
rect 213913 107883 213979 107886
rect 252369 107883 252435 107886
rect 327206 107810 327212 107812
rect 321908 107750 327212 107810
rect 327206 107748 327212 107750
rect 327276 107748 327282 107812
rect 306005 107674 306071 107677
rect 307477 107674 307543 107677
rect 306005 107672 307543 107674
rect 306005 107616 306010 107672
rect 306066 107616 307482 107672
rect 307538 107616 307543 107672
rect 306005 107614 307543 107616
rect 306005 107611 306071 107614
rect 307477 107611 307543 107614
rect 307661 107674 307727 107677
rect 307661 107672 310040 107674
rect 307661 107616 307666 107672
rect 307722 107616 310040 107672
rect 307661 107614 310040 107616
rect 307661 107611 307727 107614
rect 252461 107538 252527 107541
rect 248952 107536 252527 107538
rect 213913 106994 213979 106997
rect 217182 106994 217242 107508
rect 248952 107480 252466 107536
rect 252522 107480 252527 107536
rect 248952 107478 252527 107480
rect 252461 107475 252527 107478
rect 307661 107266 307727 107269
rect 307661 107264 310040 107266
rect 307661 107208 307666 107264
rect 307722 107208 310040 107264
rect 307661 107206 310040 107208
rect 307661 107203 307727 107206
rect 252277 106994 252343 106997
rect 213913 106992 217242 106994
rect 213913 106936 213918 106992
rect 213974 106936 217242 106992
rect 213913 106934 217242 106936
rect 248952 106992 252343 106994
rect 248952 106936 252282 106992
rect 252338 106936 252343 106992
rect 248952 106934 252343 106936
rect 213913 106931 213979 106934
rect 252277 106931 252343 106934
rect 214649 106314 214715 106317
rect 217182 106314 217242 106828
rect 309550 106754 310132 106814
rect 305729 106722 305795 106725
rect 309550 106722 309610 106754
rect 305729 106720 309610 106722
rect 305729 106664 305734 106720
rect 305790 106664 309610 106720
rect 305729 106662 309610 106664
rect 305729 106659 305795 106662
rect 252369 106586 252435 106589
rect 248952 106584 252435 106586
rect 248952 106528 252374 106584
rect 252430 106528 252435 106584
rect 248952 106526 252435 106528
rect 252369 106523 252435 106526
rect 307477 106450 307543 106453
rect 321878 106450 321938 107100
rect 342294 106450 342300 106452
rect 307477 106448 310040 106450
rect 307477 106392 307482 106448
rect 307538 106392 310040 106448
rect 307477 106390 310040 106392
rect 321878 106390 342300 106450
rect 307477 106387 307543 106390
rect 342294 106388 342300 106390
rect 342364 106388 342370 106452
rect 327022 106314 327028 106316
rect 214649 106312 217242 106314
rect 214649 106256 214654 106312
rect 214710 106256 217242 106312
rect 214649 106254 217242 106256
rect 321908 106254 327028 106314
rect 214649 106251 214715 106254
rect 327022 106252 327028 106254
rect 327092 106252 327098 106316
rect 214005 105770 214071 105773
rect 217182 105770 217242 106148
rect 252461 106042 252527 106045
rect 248952 106040 252527 106042
rect 248952 105984 252466 106040
rect 252522 105984 252527 106040
rect 248952 105982 252527 105984
rect 252461 105979 252527 105982
rect 307477 105906 307543 105909
rect 307477 105904 310040 105906
rect 307477 105848 307482 105904
rect 307538 105848 310040 105904
rect 307477 105846 310040 105848
rect 307477 105843 307543 105846
rect 214005 105768 217242 105770
rect 214005 105712 214010 105768
rect 214066 105712 217242 105768
rect 214005 105710 217242 105712
rect 214005 105707 214071 105710
rect 252277 105634 252343 105637
rect 248952 105632 252343 105634
rect 213913 105362 213979 105365
rect 217182 105362 217242 105604
rect 248952 105576 252282 105632
rect 252338 105576 252343 105632
rect 248952 105574 252343 105576
rect 252277 105571 252343 105574
rect 307661 105498 307727 105501
rect 307661 105496 310040 105498
rect 307661 105440 307666 105496
rect 307722 105440 310040 105496
rect 307661 105438 310040 105440
rect 307661 105435 307727 105438
rect 213913 105360 217242 105362
rect 213913 105304 213918 105360
rect 213974 105304 217242 105360
rect 213913 105302 217242 105304
rect 213913 105299 213979 105302
rect 214414 105164 214420 105228
rect 214484 105226 214490 105228
rect 214484 105166 217426 105226
rect 214484 105164 214490 105166
rect 217366 104924 217426 105166
rect 321510 105093 321570 105468
rect 252185 105090 252251 105093
rect 248952 105088 252251 105090
rect 248952 105032 252190 105088
rect 252246 105032 252251 105088
rect 248952 105030 252251 105032
rect 252185 105027 252251 105030
rect 307569 105090 307635 105093
rect 307569 105088 310040 105090
rect 307569 105032 307574 105088
rect 307630 105032 310040 105088
rect 307569 105030 310040 105032
rect 321510 105088 321619 105093
rect 321510 105032 321558 105088
rect 321614 105032 321619 105088
rect 321510 105030 321619 105032
rect 307569 105027 307635 105030
rect 321553 105027 321619 105030
rect 324313 104818 324379 104821
rect 321908 104816 324379 104818
rect 321908 104760 324318 104816
rect 324374 104760 324379 104816
rect 321908 104758 324379 104760
rect 324313 104755 324379 104758
rect 252461 104682 252527 104685
rect 248952 104680 252527 104682
rect 248952 104624 252466 104680
rect 252522 104624 252527 104680
rect 248952 104622 252527 104624
rect 252461 104619 252527 104622
rect 307569 104682 307635 104685
rect 307569 104680 310040 104682
rect 307569 104624 307574 104680
rect 307630 104624 310040 104680
rect 307569 104622 310040 104624
rect 307569 104619 307635 104622
rect 213913 104002 213979 104005
rect 217182 104002 217242 104244
rect 309550 104170 310132 104230
rect 252277 104138 252343 104141
rect 248952 104136 252343 104138
rect 248952 104080 252282 104136
rect 252338 104080 252343 104136
rect 248952 104078 252343 104080
rect 252277 104075 252343 104078
rect 304206 104076 304212 104140
rect 304276 104138 304282 104140
rect 309550 104138 309610 104170
rect 304276 104078 309610 104138
rect 304276 104076 304282 104078
rect 213913 104000 217242 104002
rect 213913 103944 213918 104000
rect 213974 103944 217242 104000
rect 213913 103942 217242 103944
rect 213913 103939 213979 103942
rect 307661 103866 307727 103869
rect 307661 103864 310040 103866
rect 307661 103808 307666 103864
rect 307722 103808 310040 103864
rect 307661 103806 310040 103808
rect 307661 103803 307727 103806
rect 321694 103733 321754 103972
rect 213913 103730 213979 103733
rect 252001 103730 252067 103733
rect 213913 103728 217242 103730
rect 213913 103672 213918 103728
rect 213974 103672 217242 103728
rect 213913 103670 217242 103672
rect 248952 103728 252067 103730
rect 248952 103672 252006 103728
rect 252062 103672 252067 103728
rect 248952 103670 252067 103672
rect 213913 103667 213979 103670
rect 217182 103564 217242 103670
rect 252001 103667 252067 103670
rect 321645 103728 321754 103733
rect 321645 103672 321650 103728
rect 321706 103672 321754 103728
rect 321645 103670 321754 103672
rect 321645 103667 321711 103670
rect 307569 103458 307635 103461
rect 307569 103456 310040 103458
rect 307569 103400 307574 103456
rect 307630 103400 310040 103456
rect 307569 103398 310040 103400
rect 307569 103395 307635 103398
rect 251173 103186 251239 103189
rect 323025 103186 323091 103189
rect 248952 103184 251239 103186
rect 248952 103128 251178 103184
rect 251234 103128 251239 103184
rect 248952 103126 251239 103128
rect 321908 103184 323091 103186
rect 321908 103128 323030 103184
rect 323086 103128 323091 103184
rect 321908 103126 323091 103128
rect 251173 103123 251239 103126
rect 323025 103123 323091 103126
rect 306925 103050 306991 103053
rect 306925 103048 310040 103050
rect 306925 102992 306930 103048
rect 306986 102992 310040 103048
rect 306925 102990 310040 102992
rect 306925 102987 306991 102990
rect 216213 102506 216279 102509
rect 217182 102506 217242 102884
rect 252369 102778 252435 102781
rect 248952 102776 252435 102778
rect 248952 102720 252374 102776
rect 252430 102720 252435 102776
rect 248952 102718 252435 102720
rect 252369 102715 252435 102718
rect 216213 102504 217242 102506
rect 216213 102448 216218 102504
rect 216274 102448 217242 102504
rect 216213 102446 217242 102448
rect 307661 102506 307727 102509
rect 324405 102506 324471 102509
rect 307661 102504 310040 102506
rect 307661 102448 307666 102504
rect 307722 102448 310040 102504
rect 307661 102446 310040 102448
rect 321908 102504 324471 102506
rect 321908 102448 324410 102504
rect 324466 102448 324471 102504
rect 321908 102446 324471 102448
rect 216213 102443 216279 102446
rect 307661 102443 307727 102446
rect 324405 102443 324471 102446
rect 67357 102370 67423 102373
rect 68142 102370 68816 102376
rect 67357 102368 68816 102370
rect 67357 102312 67362 102368
rect 67418 102316 68816 102368
rect 67418 102312 68202 102316
rect 67357 102310 68202 102312
rect 200070 102310 217242 102370
rect 67357 102307 67423 102310
rect 170438 102172 170444 102236
rect 170508 102234 170514 102236
rect 200070 102234 200130 102310
rect 170508 102174 200130 102234
rect 217182 102204 217242 102310
rect 252461 102234 252527 102237
rect 248952 102232 252527 102234
rect 248952 102176 252466 102232
rect 252522 102176 252527 102232
rect 248952 102174 252527 102176
rect 170508 102172 170514 102174
rect 252461 102171 252527 102174
rect 309550 101994 310132 102054
rect 304390 101900 304396 101964
rect 304460 101962 304466 101964
rect 309550 101962 309610 101994
rect 304460 101902 309610 101962
rect 304460 101900 304466 101902
rect 251357 101826 251423 101829
rect 248952 101824 251423 101826
rect 248952 101768 251362 101824
rect 251418 101768 251423 101824
rect 248952 101766 251423 101768
rect 251357 101763 251423 101766
rect 307477 101690 307543 101693
rect 307477 101688 310040 101690
rect 307477 101632 307482 101688
rect 307538 101632 310040 101688
rect 307477 101630 310040 101632
rect 307477 101627 307543 101630
rect 214557 101146 214623 101149
rect 217182 101146 217242 101524
rect 252461 101418 252527 101421
rect 248952 101416 252527 101418
rect 248952 101360 252466 101416
rect 252522 101360 252527 101416
rect 248952 101358 252527 101360
rect 252461 101355 252527 101358
rect 307569 101282 307635 101285
rect 307569 101280 310040 101282
rect 307569 101224 307574 101280
rect 307630 101224 310040 101280
rect 307569 101222 310040 101224
rect 307569 101219 307635 101222
rect 214557 101144 217242 101146
rect 214557 101088 214562 101144
rect 214618 101088 217242 101144
rect 214557 101086 217242 101088
rect 214557 101083 214623 101086
rect 321878 101010 321938 101660
rect 334014 101010 334020 101012
rect 216121 100874 216187 100877
rect 216121 100872 216874 100874
rect 216121 100816 216126 100872
rect 216182 100816 216874 100872
rect 216121 100814 216874 100816
rect 216121 100811 216187 100814
rect 67633 100738 67699 100741
rect 68142 100738 68816 100744
rect 67633 100736 68816 100738
rect 67633 100680 67638 100736
rect 67694 100684 68816 100736
rect 216814 100738 216874 100814
rect 217366 100738 217426 100980
rect 321878 100950 334020 101010
rect 334014 100948 334020 100950
rect 334084 100948 334090 101012
rect 252185 100874 252251 100877
rect 248952 100872 252251 100874
rect 248952 100816 252190 100872
rect 252246 100816 252251 100872
rect 248952 100814 252251 100816
rect 252185 100811 252251 100814
rect 307661 100874 307727 100877
rect 324262 100874 324268 100876
rect 307661 100872 310040 100874
rect 307661 100816 307666 100872
rect 307722 100816 310040 100872
rect 307661 100814 310040 100816
rect 321908 100814 324268 100874
rect 307661 100811 307727 100814
rect 324262 100812 324268 100814
rect 324332 100812 324338 100876
rect 67694 100680 68202 100684
rect 67633 100678 68202 100680
rect 216814 100678 217426 100738
rect 67633 100675 67699 100678
rect 252277 100466 252343 100469
rect 248952 100464 252343 100466
rect 248952 100408 252282 100464
rect 252338 100408 252343 100464
rect 248952 100406 252343 100408
rect 252277 100403 252343 100406
rect 307569 100466 307635 100469
rect 307569 100464 310040 100466
rect 307569 100408 307574 100464
rect 307630 100408 310040 100464
rect 307569 100406 310040 100408
rect 307569 100403 307635 100406
rect 214005 99786 214071 99789
rect 217182 99786 217242 100300
rect 324313 100194 324379 100197
rect 321908 100192 324379 100194
rect 321908 100136 324318 100192
rect 324374 100136 324379 100192
rect 321908 100134 324379 100136
rect 324313 100131 324379 100134
rect 307661 100058 307727 100061
rect 307661 100056 310040 100058
rect 307661 100000 307666 100056
rect 307722 100000 310040 100056
rect 307661 99998 310040 100000
rect 307661 99995 307727 99998
rect 252461 99922 252527 99925
rect 248952 99920 252527 99922
rect 248952 99864 252466 99920
rect 252522 99864 252527 99920
rect 248952 99862 252527 99864
rect 252461 99859 252527 99862
rect 214005 99784 217242 99786
rect 214005 99728 214010 99784
rect 214066 99728 217242 99784
rect 214005 99726 217242 99728
rect 214005 99723 214071 99726
rect 213913 99514 213979 99517
rect 213913 99512 216874 99514
rect 213913 99456 213918 99512
rect 213974 99456 216874 99512
rect 213913 99454 216874 99456
rect 213913 99451 213979 99454
rect 216814 99378 216874 99454
rect 217366 99378 217426 99620
rect 305678 99588 305684 99652
rect 305748 99650 305754 99652
rect 305748 99590 310040 99650
rect 305748 99588 305754 99590
rect 252369 99514 252435 99517
rect 248952 99512 252435 99514
rect 248952 99456 252374 99512
rect 252430 99456 252435 99512
rect 248952 99454 252435 99456
rect 252369 99451 252435 99454
rect 340086 99452 340092 99516
rect 340156 99514 340162 99516
rect 583520 99514 584960 99604
rect 340156 99454 584960 99514
rect 340156 99452 340162 99454
rect 216814 99318 217426 99378
rect 583520 99364 584960 99454
rect 307569 99106 307635 99109
rect 307569 99104 310040 99106
rect 307569 99048 307574 99104
rect 307630 99048 310040 99104
rect 307569 99046 310040 99048
rect 307569 99043 307635 99046
rect 252461 98970 252527 98973
rect 248952 98968 252527 98970
rect 214005 98426 214071 98429
rect 217182 98426 217242 98940
rect 248952 98912 252466 98968
rect 252522 98912 252527 98968
rect 248952 98910 252527 98912
rect 252461 98907 252527 98910
rect 321277 98834 321343 98837
rect 321510 98834 321570 99348
rect 321277 98832 321570 98834
rect 321277 98776 321282 98832
rect 321338 98776 321570 98832
rect 321277 98774 321570 98776
rect 321277 98771 321343 98774
rect 307017 98698 307083 98701
rect 307017 98696 310040 98698
rect 307017 98640 307022 98696
rect 307078 98640 310040 98696
rect 307017 98638 310040 98640
rect 307017 98635 307083 98638
rect 251265 98562 251331 98565
rect 248952 98560 251331 98562
rect 248952 98504 251270 98560
rect 251326 98504 251331 98560
rect 248952 98502 251331 98504
rect 251265 98499 251331 98502
rect 214005 98424 217242 98426
rect 214005 98368 214010 98424
rect 214066 98368 217242 98424
rect 214005 98366 217242 98368
rect 214005 98363 214071 98366
rect 307661 98290 307727 98293
rect 307661 98288 310040 98290
rect 166901 98020 166967 98021
rect 166901 98016 166948 98020
rect 167012 98018 167018 98020
rect 213913 98018 213979 98021
rect 217366 98018 217426 98260
rect 307661 98232 307666 98288
rect 307722 98232 310040 98288
rect 307661 98230 310040 98232
rect 307661 98227 307727 98230
rect 321878 98154 321938 98532
rect 331254 98154 331260 98156
rect 321878 98094 331260 98154
rect 331254 98092 331260 98094
rect 331324 98092 331330 98156
rect 252369 98018 252435 98021
rect 166901 97960 166906 98016
rect 166901 97956 166948 97960
rect 167012 97958 167058 98018
rect 213913 98016 217426 98018
rect 213913 97960 213918 98016
rect 213974 97960 217426 98016
rect 213913 97958 217426 97960
rect 248952 98016 252435 98018
rect 248952 97960 252374 98016
rect 252430 97960 252435 98016
rect 248952 97958 252435 97960
rect 167012 97956 167018 97958
rect 166901 97955 166967 97956
rect 213913 97955 213979 97958
rect 252369 97955 252435 97958
rect 309550 97778 310132 97838
rect -960 97610 480 97700
rect 298686 97684 298692 97748
rect 298756 97746 298762 97748
rect 309550 97746 309610 97778
rect 298756 97686 309610 97746
rect 298756 97684 298762 97686
rect 2773 97610 2839 97613
rect 252461 97610 252527 97613
rect -960 97608 2839 97610
rect -960 97552 2778 97608
rect 2834 97552 2839 97608
rect 248952 97608 252527 97610
rect -960 97550 2839 97552
rect -960 97460 480 97550
rect 2773 97547 2839 97550
rect 166390 97140 166396 97204
rect 166460 97202 166466 97204
rect 214465 97202 214531 97205
rect 166460 97200 214531 97202
rect 166460 97144 214470 97200
rect 214526 97144 214531 97200
rect 166460 97142 214531 97144
rect 166460 97140 166466 97142
rect 214465 97139 214531 97142
rect 213913 97066 213979 97069
rect 217182 97066 217242 97580
rect 248952 97552 252466 97608
rect 252522 97552 252527 97608
rect 248952 97550 252527 97552
rect 252461 97547 252527 97550
rect 307661 97474 307727 97477
rect 307661 97472 310040 97474
rect 307661 97416 307666 97472
rect 307722 97416 310040 97472
rect 307661 97414 310040 97416
rect 307661 97411 307727 97414
rect 321369 97338 321435 97341
rect 321510 97338 321570 97852
rect 321369 97336 321570 97338
rect 321369 97280 321374 97336
rect 321430 97280 321570 97336
rect 321369 97278 321570 97280
rect 321369 97275 321435 97278
rect 251265 97066 251331 97069
rect 252461 97066 252527 97069
rect 213913 97064 217242 97066
rect 213913 97008 213918 97064
rect 213974 97008 217242 97064
rect 213913 97006 217242 97008
rect 248952 97064 252527 97066
rect 248952 97008 251270 97064
rect 251326 97008 252466 97064
rect 252522 97008 252527 97064
rect 248952 97006 252527 97008
rect 213913 97003 213979 97006
rect 251265 97003 251331 97006
rect 252461 97003 252527 97006
rect 306966 97004 306972 97068
rect 307036 97066 307042 97068
rect 324497 97066 324563 97069
rect 307036 97006 310040 97066
rect 321908 97064 324563 97066
rect 321908 97008 324502 97064
rect 324558 97008 324563 97064
rect 321908 97006 324563 97008
rect 307036 97004 307042 97006
rect 324497 97003 324563 97006
rect 214925 96658 214991 96661
rect 217182 96658 217242 96900
rect 262806 96794 262812 96796
rect 251958 96734 262812 96794
rect 249149 96658 249215 96661
rect 251958 96658 252018 96734
rect 262806 96732 262812 96734
rect 262876 96732 262882 96796
rect 214925 96656 217242 96658
rect 214925 96600 214930 96656
rect 214986 96600 217242 96656
rect 214925 96598 217242 96600
rect 248952 96656 252018 96658
rect 248952 96600 249154 96656
rect 249210 96600 252018 96656
rect 248952 96598 252018 96600
rect 252461 96658 252527 96661
rect 260046 96658 260052 96660
rect 252461 96656 260052 96658
rect 252461 96600 252466 96656
rect 252522 96600 260052 96656
rect 252461 96598 260052 96600
rect 214925 96595 214991 96598
rect 249149 96595 249215 96598
rect 252461 96595 252527 96598
rect 260046 96596 260052 96598
rect 260116 96596 260122 96660
rect 306925 96658 306991 96661
rect 321461 96658 321527 96661
rect 306925 96656 310040 96658
rect 306925 96600 306930 96656
rect 306986 96600 310040 96656
rect 306925 96598 310040 96600
rect 321461 96656 321570 96658
rect 321461 96600 321466 96656
rect 321522 96600 321570 96656
rect 306925 96595 306991 96598
rect 321461 96595 321570 96600
rect 321510 96356 321570 96595
rect 213913 95842 213979 95845
rect 217182 95842 217242 96356
rect 251173 96250 251239 96253
rect 248860 96248 251239 96250
rect 248860 96192 251178 96248
rect 251234 96192 251239 96248
rect 248860 96190 251239 96192
rect 251173 96187 251239 96190
rect 307661 96250 307727 96253
rect 307661 96248 310132 96250
rect 307661 96192 307666 96248
rect 307722 96192 310132 96248
rect 307661 96190 310132 96192
rect 307661 96187 307727 96190
rect 213913 95840 217242 95842
rect 213913 95784 213918 95840
rect 213974 95784 217242 95840
rect 213913 95782 217242 95784
rect 213913 95779 213979 95782
rect 164877 95162 164943 95165
rect 166942 95162 166948 95164
rect 164877 95160 166948 95162
rect 164877 95104 164882 95160
rect 164938 95104 166948 95160
rect 164877 95102 166948 95104
rect 164877 95099 164943 95102
rect 166942 95100 166948 95102
rect 167012 95100 167018 95164
rect 177297 95162 177363 95165
rect 321277 95162 321343 95165
rect 177297 95160 321343 95162
rect 177297 95104 177302 95160
rect 177358 95104 321282 95160
rect 321338 95104 321343 95160
rect 177297 95102 321343 95104
rect 177297 95099 177363 95102
rect 321277 95099 321343 95102
rect 66161 94890 66227 94893
rect 207749 94890 207815 94893
rect 66161 94888 207815 94890
rect 66161 94832 66166 94888
rect 66222 94832 207754 94888
rect 207810 94832 207815 94888
rect 66161 94830 207815 94832
rect 66161 94827 66227 94830
rect 207749 94827 207815 94830
rect 111977 94756 112043 94757
rect 113725 94756 113791 94757
rect 129365 94756 129431 94757
rect 151629 94756 151695 94757
rect 111912 94692 111918 94756
rect 111982 94754 112043 94756
rect 111982 94752 112074 94754
rect 112038 94696 112074 94752
rect 111982 94694 112074 94696
rect 111982 94692 112043 94694
rect 113680 94692 113686 94756
rect 113750 94754 113791 94756
rect 113750 94752 113842 94754
rect 113786 94696 113842 94752
rect 113750 94694 113842 94696
rect 113750 94692 113791 94694
rect 129320 94692 129326 94756
rect 129390 94754 129431 94756
rect 151624 94754 151630 94756
rect 129390 94752 129482 94754
rect 129426 94696 129482 94752
rect 129390 94694 129482 94696
rect 151538 94694 151630 94754
rect 129390 94692 129431 94694
rect 151624 94692 151630 94694
rect 151694 94692 151700 94756
rect 111977 94691 112043 94692
rect 113725 94691 113791 94692
rect 129365 94691 129431 94692
rect 151629 94691 151695 94692
rect 161473 94482 161539 94485
rect 199377 94482 199443 94485
rect 161473 94480 199443 94482
rect 161473 94424 161478 94480
rect 161534 94424 199382 94480
rect 199438 94424 199443 94480
rect 161473 94422 199443 94424
rect 161473 94419 161539 94422
rect 199377 94419 199443 94422
rect 67541 93802 67607 93805
rect 214414 93802 214420 93804
rect 67541 93800 214420 93802
rect 67541 93744 67546 93800
rect 67602 93744 214420 93800
rect 67541 93742 214420 93744
rect 67541 93739 67607 93742
rect 214414 93740 214420 93742
rect 214484 93740 214490 93804
rect 118049 93668 118115 93669
rect 133137 93668 133203 93669
rect 117998 93666 118004 93668
rect 117958 93606 118004 93666
rect 118068 93664 118115 93668
rect 133086 93666 133092 93668
rect 118110 93608 118115 93664
rect 117998 93604 118004 93606
rect 118068 93604 118115 93608
rect 133046 93606 133092 93666
rect 133156 93664 133203 93668
rect 133198 93608 133203 93664
rect 133086 93604 133092 93606
rect 133156 93604 133203 93608
rect 118049 93603 118115 93604
rect 133137 93603 133203 93604
rect 85665 93532 85731 93533
rect 107745 93532 107811 93533
rect 120625 93532 120691 93533
rect 85614 93530 85620 93532
rect 85574 93470 85620 93530
rect 85684 93528 85731 93532
rect 107694 93530 107700 93532
rect 85726 93472 85731 93528
rect 85614 93468 85620 93470
rect 85684 93468 85731 93472
rect 107654 93470 107700 93530
rect 107764 93528 107811 93532
rect 120574 93530 120580 93532
rect 107806 93472 107811 93528
rect 107694 93468 107700 93470
rect 107764 93468 107811 93472
rect 120534 93470 120580 93530
rect 120644 93528 120691 93532
rect 120686 93472 120691 93528
rect 120574 93468 120580 93470
rect 120644 93468 120691 93472
rect 85665 93467 85731 93468
rect 107745 93467 107811 93468
rect 120625 93467 120691 93468
rect 110137 93260 110203 93261
rect 110086 93258 110092 93260
rect 110046 93198 110092 93258
rect 110156 93256 110203 93260
rect 110198 93200 110203 93256
rect 110086 93196 110092 93198
rect 110156 93196 110203 93200
rect 110137 93195 110203 93196
rect 84326 92380 84332 92444
rect 84396 92442 84402 92444
rect 85113 92442 85179 92445
rect 84396 92440 85179 92442
rect 84396 92384 85118 92440
rect 85174 92384 85179 92440
rect 84396 92382 85179 92384
rect 84396 92380 84402 92382
rect 85113 92379 85179 92382
rect 91318 92380 91324 92444
rect 91388 92442 91394 92444
rect 91645 92442 91711 92445
rect 95049 92444 95115 92445
rect 94998 92442 95004 92444
rect 91388 92440 91711 92442
rect 91388 92384 91650 92440
rect 91706 92384 91711 92440
rect 91388 92382 91711 92384
rect 94958 92382 95004 92442
rect 95068 92440 95115 92444
rect 95110 92384 95115 92440
rect 91388 92380 91394 92382
rect 91645 92379 91711 92382
rect 94998 92380 95004 92382
rect 95068 92380 95115 92384
rect 105670 92380 105676 92444
rect 105740 92442 105746 92444
rect 105997 92442 106063 92445
rect 115473 92444 115539 92445
rect 116761 92444 116827 92445
rect 115422 92442 115428 92444
rect 105740 92440 106063 92442
rect 105740 92384 106002 92440
rect 106058 92384 106063 92440
rect 105740 92382 106063 92384
rect 115382 92382 115428 92442
rect 115492 92440 115539 92444
rect 116710 92442 116716 92444
rect 115534 92384 115539 92440
rect 105740 92380 105746 92382
rect 95049 92379 95115 92380
rect 105997 92379 106063 92382
rect 115422 92380 115428 92382
rect 115492 92380 115539 92384
rect 116670 92382 116716 92442
rect 116780 92440 116827 92444
rect 116822 92384 116827 92440
rect 116710 92380 116716 92382
rect 116780 92380 116827 92384
rect 120206 92380 120212 92444
rect 120276 92442 120282 92444
rect 120533 92442 120599 92445
rect 120276 92440 120599 92442
rect 120276 92384 120538 92440
rect 120594 92384 120599 92440
rect 120276 92382 120599 92384
rect 120276 92380 120282 92382
rect 115473 92379 115539 92380
rect 116761 92379 116827 92380
rect 120533 92379 120599 92382
rect 125358 92380 125364 92444
rect 125428 92442 125434 92444
rect 125501 92442 125567 92445
rect 125961 92444 126027 92445
rect 130745 92444 130811 92445
rect 151721 92444 151787 92445
rect 152089 92444 152155 92445
rect 125910 92442 125916 92444
rect 125428 92440 125567 92442
rect 125428 92384 125506 92440
rect 125562 92384 125567 92440
rect 125428 92382 125567 92384
rect 125870 92382 125916 92442
rect 125980 92440 126027 92444
rect 130694 92442 130700 92444
rect 126022 92384 126027 92440
rect 125428 92380 125434 92382
rect 125501 92379 125567 92382
rect 125910 92380 125916 92382
rect 125980 92380 126027 92384
rect 130654 92382 130700 92442
rect 130764 92440 130811 92444
rect 151670 92442 151676 92444
rect 130806 92384 130811 92440
rect 130694 92380 130700 92382
rect 130764 92380 130811 92384
rect 151630 92382 151676 92442
rect 151740 92440 151787 92444
rect 152038 92442 152044 92444
rect 151782 92384 151787 92440
rect 151670 92380 151676 92382
rect 151740 92380 151787 92384
rect 151998 92382 152044 92442
rect 152108 92440 152155 92444
rect 152150 92384 152155 92440
rect 152038 92380 152044 92382
rect 152108 92380 152155 92384
rect 125961 92379 126027 92380
rect 130745 92379 130811 92380
rect 151721 92379 151787 92380
rect 152089 92379 152155 92380
rect 109166 92244 109172 92308
rect 109236 92306 109242 92308
rect 110321 92306 110387 92309
rect 109236 92304 110387 92306
rect 109236 92248 110326 92304
rect 110382 92248 110387 92304
rect 109236 92246 110387 92248
rect 109236 92244 109242 92246
rect 110321 92243 110387 92246
rect 119286 92244 119292 92308
rect 119356 92306 119362 92308
rect 166390 92306 166396 92308
rect 119356 92246 166396 92306
rect 119356 92244 119362 92246
rect 166390 92244 166396 92246
rect 166460 92244 166466 92308
rect 136030 92108 136036 92172
rect 136100 92170 136106 92172
rect 136449 92170 136515 92173
rect 136100 92168 136515 92170
rect 136100 92112 136454 92168
rect 136510 92112 136515 92168
rect 136100 92110 136515 92112
rect 136100 92108 136106 92110
rect 136449 92107 136515 92110
rect 90214 91700 90220 91764
rect 90284 91762 90290 91764
rect 90633 91762 90699 91765
rect 90284 91760 90699 91762
rect 90284 91704 90638 91760
rect 90694 91704 90699 91760
rect 90284 91702 90699 91704
rect 90284 91700 90290 91702
rect 90633 91699 90699 91702
rect 102542 91700 102548 91764
rect 102612 91762 102618 91764
rect 102685 91762 102751 91765
rect 102612 91760 102751 91762
rect 102612 91704 102690 91760
rect 102746 91704 102751 91760
rect 102612 91702 102751 91704
rect 102612 91700 102618 91702
rect 102685 91699 102751 91702
rect 114870 91700 114876 91764
rect 114940 91762 114946 91764
rect 115381 91762 115447 91765
rect 126697 91764 126763 91765
rect 126646 91762 126652 91764
rect 114940 91760 115447 91762
rect 114940 91704 115386 91760
rect 115442 91704 115447 91760
rect 114940 91702 115447 91704
rect 126606 91702 126652 91762
rect 126716 91760 126763 91764
rect 126758 91704 126763 91760
rect 114940 91700 114946 91702
rect 115381 91699 115447 91702
rect 126646 91700 126652 91702
rect 126716 91700 126763 91704
rect 126697 91699 126763 91700
rect 100017 91628 100083 91629
rect 99966 91626 99972 91628
rect 99926 91566 99972 91626
rect 100036 91624 100083 91628
rect 100078 91568 100083 91624
rect 99966 91564 99972 91566
rect 100036 91564 100083 91568
rect 102726 91564 102732 91628
rect 102796 91626 102802 91628
rect 161473 91626 161539 91629
rect 102796 91624 161539 91626
rect 102796 91568 161478 91624
rect 161534 91568 161539 91624
rect 102796 91566 161539 91568
rect 102796 91564 102802 91566
rect 100017 91563 100083 91564
rect 161473 91563 161539 91566
rect 98126 91428 98132 91492
rect 98196 91490 98202 91492
rect 99281 91490 99347 91493
rect 101857 91492 101923 91493
rect 122833 91492 122899 91493
rect 101806 91490 101812 91492
rect 98196 91488 99347 91490
rect 98196 91432 99286 91488
rect 99342 91432 99347 91488
rect 98196 91430 99347 91432
rect 101766 91430 101812 91490
rect 101876 91488 101923 91492
rect 101918 91432 101923 91488
rect 98196 91428 98202 91430
rect 99281 91427 99347 91430
rect 101806 91428 101812 91430
rect 101876 91428 101923 91432
rect 122782 91428 122788 91492
rect 122852 91490 122899 91492
rect 122852 91488 122944 91490
rect 122894 91432 122944 91488
rect 122852 91430 122944 91432
rect 122852 91428 122899 91430
rect 151118 91428 151124 91492
rect 151188 91490 151194 91492
rect 151261 91490 151327 91493
rect 151188 91488 151327 91490
rect 151188 91432 151266 91488
rect 151322 91432 151327 91488
rect 151188 91430 151327 91432
rect 151188 91428 151194 91430
rect 101857 91427 101923 91428
rect 122833 91427 122899 91428
rect 151261 91427 151327 91430
rect 96654 91292 96660 91356
rect 96724 91354 96730 91356
rect 97809 91354 97875 91357
rect 96724 91352 97875 91354
rect 96724 91296 97814 91352
rect 97870 91296 97875 91352
rect 96724 91294 97875 91296
rect 96724 91292 96730 91294
rect 97809 91291 97875 91294
rect 98494 91292 98500 91356
rect 98564 91354 98570 91356
rect 99097 91354 99163 91357
rect 98564 91352 99163 91354
rect 98564 91296 99102 91352
rect 99158 91296 99163 91352
rect 98564 91294 99163 91296
rect 98564 91292 98570 91294
rect 99097 91291 99163 91294
rect 100886 91292 100892 91356
rect 100956 91354 100962 91356
rect 102041 91354 102107 91357
rect 100956 91352 102107 91354
rect 100956 91296 102046 91352
rect 102102 91296 102107 91352
rect 100956 91294 102107 91296
rect 100956 91292 100962 91294
rect 102041 91291 102107 91294
rect 106406 91292 106412 91356
rect 106476 91354 106482 91356
rect 107561 91354 107627 91357
rect 106476 91352 107627 91354
rect 106476 91296 107566 91352
rect 107622 91296 107627 91352
rect 106476 91294 107627 91296
rect 106476 91292 106482 91294
rect 107561 91291 107627 91294
rect 111190 91292 111196 91356
rect 111260 91354 111266 91356
rect 111425 91354 111491 91357
rect 114369 91356 114435 91357
rect 114318 91354 114324 91356
rect 111260 91352 111491 91354
rect 111260 91296 111430 91352
rect 111486 91296 111491 91352
rect 111260 91294 111491 91296
rect 114278 91294 114324 91354
rect 114388 91352 114435 91356
rect 114430 91296 114435 91352
rect 111260 91292 111266 91294
rect 111425 91291 111491 91294
rect 114318 91292 114324 91294
rect 114388 91292 114435 91296
rect 121678 91292 121684 91356
rect 121748 91354 121754 91356
rect 122741 91354 122807 91357
rect 121748 91352 122807 91354
rect 121748 91296 122746 91352
rect 122802 91296 122807 91352
rect 121748 91294 122807 91296
rect 121748 91292 121754 91294
rect 114369 91291 114435 91292
rect 122741 91291 122807 91294
rect 74758 91156 74764 91220
rect 74828 91218 74834 91220
rect 75821 91218 75887 91221
rect 74828 91216 75887 91218
rect 74828 91160 75826 91216
rect 75882 91160 75887 91216
rect 74828 91158 75887 91160
rect 74828 91156 74834 91158
rect 75821 91155 75887 91158
rect 86718 91156 86724 91220
rect 86788 91218 86794 91220
rect 86861 91218 86927 91221
rect 88057 91220 88123 91221
rect 88006 91218 88012 91220
rect 86788 91216 86927 91218
rect 86788 91160 86866 91216
rect 86922 91160 86927 91216
rect 86788 91158 86927 91160
rect 87966 91158 88012 91218
rect 88076 91216 88123 91220
rect 88118 91160 88123 91216
rect 86788 91156 86794 91158
rect 86861 91155 86927 91158
rect 88006 91156 88012 91158
rect 88076 91156 88123 91160
rect 88926 91156 88932 91220
rect 88996 91218 89002 91220
rect 89621 91218 89687 91221
rect 88996 91216 89687 91218
rect 88996 91160 89626 91216
rect 89682 91160 89687 91216
rect 88996 91158 89687 91160
rect 88996 91156 89002 91158
rect 88057 91155 88123 91156
rect 89621 91155 89687 91158
rect 92606 91156 92612 91220
rect 92676 91218 92682 91220
rect 93761 91218 93827 91221
rect 92676 91216 93827 91218
rect 92676 91160 93766 91216
rect 93822 91160 93827 91216
rect 92676 91158 93827 91160
rect 92676 91156 92682 91158
rect 93761 91155 93827 91158
rect 93894 91156 93900 91220
rect 93964 91218 93970 91220
rect 95141 91218 95207 91221
rect 93964 91216 95207 91218
rect 93964 91160 95146 91216
rect 95202 91160 95207 91216
rect 93964 91158 95207 91160
rect 93964 91156 93970 91158
rect 95141 91155 95207 91158
rect 96286 91156 96292 91220
rect 96356 91218 96362 91220
rect 96521 91218 96587 91221
rect 96356 91216 96587 91218
rect 96356 91160 96526 91216
rect 96582 91160 96587 91216
rect 96356 91158 96587 91160
rect 96356 91156 96362 91158
rect 96521 91155 96587 91158
rect 97206 91156 97212 91220
rect 97276 91218 97282 91220
rect 97901 91218 97967 91221
rect 97276 91216 97967 91218
rect 97276 91160 97906 91216
rect 97962 91160 97967 91216
rect 97276 91158 97967 91160
rect 97276 91156 97282 91158
rect 97901 91155 97967 91158
rect 99046 91156 99052 91220
rect 99116 91218 99122 91220
rect 99189 91218 99255 91221
rect 100569 91220 100635 91221
rect 100518 91218 100524 91220
rect 99116 91216 99255 91218
rect 99116 91160 99194 91216
rect 99250 91160 99255 91216
rect 99116 91158 99255 91160
rect 100478 91158 100524 91218
rect 100588 91216 100635 91220
rect 101949 91220 102015 91221
rect 104249 91220 104315 91221
rect 101949 91218 101996 91220
rect 100630 91160 100635 91216
rect 99116 91156 99122 91158
rect 99189 91155 99255 91158
rect 100518 91156 100524 91158
rect 100588 91156 100635 91160
rect 101904 91216 101996 91218
rect 101904 91160 101954 91216
rect 101904 91158 101996 91160
rect 100569 91155 100635 91156
rect 101949 91156 101996 91158
rect 102060 91156 102066 91220
rect 104198 91218 104204 91220
rect 104158 91158 104204 91218
rect 104268 91216 104315 91220
rect 104310 91160 104315 91216
rect 104198 91156 104204 91158
rect 104268 91156 104315 91160
rect 104566 91156 104572 91220
rect 104636 91218 104642 91220
rect 104801 91218 104867 91221
rect 104636 91216 104867 91218
rect 104636 91160 104806 91216
rect 104862 91160 104867 91216
rect 104636 91158 104867 91160
rect 104636 91156 104642 91158
rect 101949 91155 102015 91156
rect 104249 91155 104315 91156
rect 104801 91155 104867 91158
rect 105486 91156 105492 91220
rect 105556 91218 105562 91220
rect 106181 91218 106247 91221
rect 105556 91216 106247 91218
rect 105556 91160 106186 91216
rect 106242 91160 106247 91216
rect 105556 91158 106247 91160
rect 105556 91156 105562 91158
rect 106181 91155 106247 91158
rect 106774 91156 106780 91220
rect 106844 91218 106850 91220
rect 107469 91218 107535 91221
rect 106844 91216 107535 91218
rect 106844 91160 107474 91216
rect 107530 91160 107535 91216
rect 106844 91158 107535 91160
rect 106844 91156 106850 91158
rect 107469 91155 107535 91158
rect 108062 91156 108068 91220
rect 108132 91218 108138 91220
rect 108941 91218 109007 91221
rect 109585 91220 109651 91221
rect 109534 91218 109540 91220
rect 108132 91216 109007 91218
rect 108132 91160 108946 91216
rect 109002 91160 109007 91216
rect 108132 91158 109007 91160
rect 109494 91158 109540 91218
rect 109604 91216 109651 91220
rect 109646 91160 109651 91216
rect 108132 91156 108138 91158
rect 108941 91155 109007 91158
rect 109534 91156 109540 91158
rect 109604 91156 109651 91160
rect 110638 91156 110644 91220
rect 110708 91218 110714 91220
rect 111241 91218 111307 91221
rect 112345 91220 112411 91221
rect 112294 91218 112300 91220
rect 110708 91216 111307 91218
rect 110708 91160 111246 91216
rect 111302 91160 111307 91216
rect 110708 91158 111307 91160
rect 112254 91158 112300 91218
rect 112364 91216 112411 91220
rect 112406 91160 112411 91216
rect 110708 91156 110714 91158
rect 109585 91155 109651 91156
rect 111241 91155 111307 91158
rect 112294 91156 112300 91158
rect 112364 91156 112411 91160
rect 113214 91156 113220 91220
rect 113284 91218 113290 91220
rect 114461 91218 114527 91221
rect 115841 91220 115907 91221
rect 117129 91220 117195 91221
rect 115790 91218 115796 91220
rect 113284 91216 114527 91218
rect 113284 91160 114466 91216
rect 114522 91160 114527 91216
rect 113284 91158 114527 91160
rect 115750 91158 115796 91218
rect 115860 91216 115907 91220
rect 117078 91218 117084 91220
rect 115902 91160 115907 91216
rect 113284 91156 113290 91158
rect 112345 91155 112411 91156
rect 114461 91155 114527 91158
rect 115790 91156 115796 91158
rect 115860 91156 115907 91160
rect 117038 91158 117084 91218
rect 117148 91216 117195 91220
rect 117190 91160 117195 91216
rect 117078 91156 117084 91158
rect 117148 91156 117195 91160
rect 118182 91156 118188 91220
rect 118252 91218 118258 91220
rect 118601 91218 118667 91221
rect 118252 91216 118667 91218
rect 118252 91160 118606 91216
rect 118662 91160 118667 91216
rect 118252 91158 118667 91160
rect 118252 91156 118258 91158
rect 115841 91155 115907 91156
rect 117129 91155 117195 91156
rect 118601 91155 118667 91158
rect 119654 91156 119660 91220
rect 119724 91218 119730 91220
rect 119981 91218 120047 91221
rect 119724 91216 120047 91218
rect 119724 91160 119986 91216
rect 120042 91160 120047 91216
rect 119724 91158 120047 91160
rect 119724 91156 119730 91158
rect 119981 91155 120047 91158
rect 122046 91156 122052 91220
rect 122116 91218 122122 91220
rect 122649 91218 122715 91221
rect 122116 91216 122715 91218
rect 122116 91160 122654 91216
rect 122710 91160 122715 91216
rect 122116 91158 122715 91160
rect 122116 91156 122122 91158
rect 122649 91155 122715 91158
rect 123150 91156 123156 91220
rect 123220 91218 123226 91220
rect 123477 91218 123543 91221
rect 124121 91220 124187 91221
rect 124070 91218 124076 91220
rect 123220 91216 123543 91218
rect 123220 91160 123482 91216
rect 123538 91160 123543 91216
rect 123220 91158 123543 91160
rect 124030 91158 124076 91218
rect 124140 91216 124187 91220
rect 124182 91160 124187 91216
rect 123220 91156 123226 91158
rect 123477 91155 123543 91158
rect 124070 91156 124076 91158
rect 124140 91156 124187 91160
rect 124438 91156 124444 91220
rect 124508 91218 124514 91220
rect 125409 91218 125475 91221
rect 126513 91220 126579 91221
rect 126462 91218 126468 91220
rect 124508 91216 125475 91218
rect 124508 91160 125414 91216
rect 125470 91160 125475 91216
rect 124508 91158 125475 91160
rect 126422 91158 126468 91218
rect 126532 91216 126579 91220
rect 126574 91160 126579 91216
rect 124508 91156 124514 91158
rect 124121 91155 124187 91156
rect 125409 91155 125475 91158
rect 126462 91156 126468 91158
rect 126532 91156 126579 91160
rect 127566 91156 127572 91220
rect 127636 91218 127642 91220
rect 128261 91218 128327 91221
rect 132401 91220 132467 91221
rect 132350 91218 132356 91220
rect 127636 91216 128327 91218
rect 127636 91160 128266 91216
rect 128322 91160 128327 91216
rect 127636 91158 128327 91160
rect 132310 91158 132356 91218
rect 132420 91216 132467 91220
rect 132462 91160 132467 91216
rect 127636 91156 127642 91158
rect 126513 91155 126579 91156
rect 128261 91155 128327 91158
rect 132350 91156 132356 91158
rect 132420 91156 132467 91160
rect 134374 91156 134380 91220
rect 134444 91218 134450 91220
rect 134609 91218 134675 91221
rect 134444 91216 134675 91218
rect 134444 91160 134614 91216
rect 134670 91160 134675 91216
rect 134444 91158 134675 91160
rect 134444 91156 134450 91158
rect 132401 91155 132467 91156
rect 134609 91155 134675 91158
rect 65977 91082 66043 91085
rect 170438 91082 170444 91084
rect 65977 91080 170444 91082
rect 65977 91024 65982 91080
rect 66038 91024 170444 91080
rect 65977 91022 170444 91024
rect 65977 91019 66043 91022
rect 170438 91020 170444 91022
rect 170508 91020 170514 91084
rect 126697 89722 126763 89725
rect 168966 89722 168972 89724
rect 126697 89720 168972 89722
rect 126697 89664 126702 89720
rect 126758 89664 168972 89720
rect 126697 89662 168972 89664
rect 126697 89659 126763 89662
rect 168966 89660 168972 89662
rect 169036 89660 169042 89724
rect 114369 88226 114435 88229
rect 166206 88226 166212 88228
rect 114369 88224 166212 88226
rect 114369 88168 114374 88224
rect 114430 88168 166212 88224
rect 114369 88166 166212 88168
rect 114369 88163 114435 88166
rect 166206 88164 166212 88166
rect 166276 88164 166282 88228
rect 582833 86186 582899 86189
rect 583520 86186 584960 86276
rect 582833 86184 584960 86186
rect 582833 86128 582838 86184
rect 582894 86128 584960 86184
rect 582833 86126 584960 86128
rect 582833 86123 582899 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 97809 81426 97875 81429
rect 173014 81426 173020 81428
rect 97809 81424 173020 81426
rect 97809 81368 97814 81424
rect 97870 81368 173020 81424
rect 97809 81366 173020 81368
rect 97809 81363 97875 81366
rect 173014 81364 173020 81366
rect 173084 81364 173090 81428
rect 99189 80066 99255 80069
rect 170254 80066 170260 80068
rect 99189 80064 170260 80066
rect 99189 80008 99194 80064
rect 99250 80008 170260 80064
rect 99189 80006 170260 80008
rect 99189 80003 99255 80006
rect 170254 80004 170260 80006
rect 170324 80004 170330 80068
rect 99281 78570 99347 78573
rect 169150 78570 169156 78572
rect 99281 78568 169156 78570
rect 99281 78512 99286 78568
rect 99342 78512 169156 78568
rect 99281 78510 169156 78512
rect 99281 78507 99347 78510
rect 169150 78508 169156 78510
rect 169220 78508 169226 78572
rect 580257 72994 580323 72997
rect 583520 72994 584960 73084
rect 580257 72992 584960 72994
rect 580257 72936 580262 72992
rect 580318 72936 584960 72992
rect 580257 72934 584960 72936
rect 580257 72931 580323 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3509 71634 3575 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 35893 62794 35959 62797
rect 304390 62794 304396 62796
rect 35893 62792 304396 62794
rect 35893 62736 35898 62792
rect 35954 62736 304396 62792
rect 35893 62734 304396 62736
rect 35893 62731 35959 62734
rect 304390 62732 304396 62734
rect 304460 62732 304466 62796
rect 8293 61434 8359 61437
rect 302918 61434 302924 61436
rect 8293 61432 302924 61434
rect 8293 61376 8298 61432
rect 8354 61376 302924 61432
rect 8293 61374 302924 61376
rect 8293 61371 8359 61374
rect 302918 61372 302924 61374
rect 302988 61372 302994 61436
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3417 58578 3483 58581
rect -960 58576 3483 58578
rect -960 58520 3422 58576
rect 3478 58520 3483 58576
rect -960 58518 3483 58520
rect -960 58428 480 58518
rect 3417 58515 3483 58518
rect 15193 57218 15259 57221
rect 298686 57218 298692 57220
rect 15193 57216 298692 57218
rect 15193 57160 15198 57216
rect 15254 57160 298692 57216
rect 15193 57158 298692 57160
rect 15193 57155 15259 57158
rect 298686 57156 298692 57158
rect 298756 57156 298762 57220
rect 12433 54498 12499 54501
rect 301814 54498 301820 54500
rect 12433 54496 301820 54498
rect 12433 54440 12438 54496
rect 12494 54440 301820 54496
rect 12433 54438 301820 54440
rect 12433 54435 12499 54438
rect 301814 54436 301820 54438
rect 301884 54436 301890 54500
rect 49693 47562 49759 47565
rect 305494 47562 305500 47564
rect 49693 47560 305500 47562
rect 49693 47504 49698 47560
rect 49754 47504 305500 47560
rect 49693 47502 305500 47504
rect 49693 47499 49759 47502
rect 305494 47500 305500 47502
rect 305564 47500 305570 47564
rect 583109 46338 583175 46341
rect 583520 46338 584960 46428
rect 583109 46336 584960 46338
rect 583109 46280 583114 46336
rect 583170 46280 584960 46336
rect 583109 46278 584960 46280
rect 583109 46275 583175 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 582557 33146 582623 33149
rect 583520 33146 584960 33236
rect 582557 33144 584960 33146
rect 582557 33088 582562 33144
rect 582618 33088 584960 33144
rect 582557 33086 584960 33088
rect 582557 33083 582623 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3141 32466 3207 32469
rect -960 32464 3207 32466
rect -960 32408 3146 32464
rect 3202 32408 3207 32464
rect -960 32406 3207 32408
rect -960 32316 480 32406
rect 3141 32403 3207 32406
rect 47577 32466 47643 32469
rect 307150 32466 307156 32468
rect 47577 32464 307156 32466
rect 47577 32408 47582 32464
rect 47638 32408 307156 32464
rect 47577 32406 307156 32408
rect 47577 32403 47643 32406
rect 307150 32404 307156 32406
rect 307220 32404 307226 32468
rect 59353 30970 59419 30973
rect 299974 30970 299980 30972
rect 59353 30968 299980 30970
rect 59353 30912 59358 30968
rect 59414 30912 299980 30968
rect 59353 30910 299980 30912
rect 59353 30907 59419 30910
rect 299974 30908 299980 30910
rect 300044 30908 300050 30972
rect 77385 29610 77451 29613
rect 302734 29610 302740 29612
rect 77385 29608 302740 29610
rect 77385 29552 77390 29608
rect 77446 29552 302740 29608
rect 77385 29550 302740 29552
rect 77385 29547 77451 29550
rect 302734 29548 302740 29550
rect 302804 29548 302810 29612
rect 582465 19818 582531 19821
rect 583520 19818 584960 19908
rect 582465 19816 584960 19818
rect 582465 19760 582470 19816
rect 582526 19760 584960 19816
rect 582465 19758 584960 19760
rect 582465 19755 582531 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 11053 18594 11119 18597
rect 305678 18594 305684 18596
rect 11053 18592 305684 18594
rect 11053 18536 11058 18592
rect 11114 18536 305684 18592
rect 11053 18534 305684 18536
rect 11053 18531 11119 18534
rect 305678 18532 305684 18534
rect 305748 18532 305754 18596
rect 54937 13018 55003 13021
rect 304206 13018 304212 13020
rect 54937 13016 304212 13018
rect 54937 12960 54942 13016
rect 54998 12960 304212 13016
rect 54937 12958 304212 12960
rect 54937 12955 55003 12958
rect 304206 12956 304212 12958
rect 304276 12956 304282 13020
rect 582373 6626 582439 6629
rect 583520 6626 584960 6716
rect 582373 6624 584960 6626
rect -960 6490 480 6580
rect 582373 6568 582378 6624
rect 582434 6568 584960 6624
rect 582373 6566 584960 6568
rect 582373 6563 582439 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 6453 4858 6519 4861
rect 306966 4858 306972 4860
rect 6453 4856 306972 4858
rect 6453 4800 6458 4856
rect 6514 4800 306972 4856
rect 6453 4798 306972 4800
rect 6453 4795 6519 4798
rect 306966 4796 306972 4798
rect 307036 4796 307042 4860
<< via3 >>
rect 70900 702476 70964 702540
rect 59124 700300 59188 700364
rect 61884 456860 61948 456924
rect 68876 313924 68940 313988
rect 331260 300868 331324 300932
rect 254532 296788 254596 296852
rect 120028 293932 120092 293996
rect 335124 291892 335188 291956
rect 342116 291212 342180 291276
rect 120028 289172 120092 289236
rect 70532 288764 70596 288828
rect 68876 288356 68940 288420
rect 122052 287676 122116 287740
rect 64644 284412 64708 284476
rect 166948 271900 167012 271964
rect 122052 269724 122116 269788
rect 263548 269180 263612 269244
rect 340092 264148 340156 264212
rect 338620 259524 338684 259588
rect 66116 256668 66180 256732
rect 62988 254084 63052 254148
rect 120028 253132 120092 253196
rect 258396 245652 258460 245716
rect 59124 241708 59188 241772
rect 61884 240348 61948 240412
rect 120028 239804 120092 239868
rect 66116 236540 66180 236604
rect 345060 236540 345124 236604
rect 62988 232460 63052 232524
rect 64644 226884 64708 226948
rect 320220 225524 320284 225588
rect 327028 222804 327092 222868
rect 267780 218588 267844 218652
rect 327212 213148 327276 213212
rect 342300 211788 342364 211852
rect 334020 210292 334084 210356
rect 269068 203492 269132 203556
rect 324268 196556 324332 196620
rect 336780 194516 336844 194580
rect 266308 192476 266372 192540
rect 263732 190980 263796 191044
rect 256740 185540 256804 185604
rect 166212 183636 166276 183700
rect 335492 179964 335556 180028
rect 166396 179420 166460 179484
rect 338252 179344 338316 179348
rect 338252 179288 338302 179344
rect 338302 179288 338316 179344
rect 338252 179284 338316 179288
rect 334204 178876 334268 178940
rect 255268 178740 255332 178804
rect 332548 178740 332612 178804
rect 97028 177652 97092 177716
rect 98316 177652 98380 177716
rect 105676 177652 105740 177716
rect 106964 177652 107028 177716
rect 114324 177652 114388 177716
rect 116900 177712 116964 177716
rect 116900 177656 116950 177712
rect 116950 177656 116964 177712
rect 116900 177652 116964 177656
rect 118372 177652 118436 177716
rect 120764 177652 120828 177716
rect 129412 177712 129476 177716
rect 129412 177656 129462 177712
rect 129462 177656 129476 177712
rect 129412 177652 129476 177656
rect 132356 177712 132420 177716
rect 132356 177656 132406 177712
rect 132406 177656 132420 177712
rect 132356 177652 132420 177656
rect 133092 177652 133156 177716
rect 258396 177516 258460 177580
rect 259500 177380 259564 177444
rect 249380 177244 249444 177308
rect 331444 177244 331508 177308
rect 112116 177108 112180 177172
rect 110644 177032 110708 177036
rect 110644 176976 110694 177032
rect 110694 176976 110708 177032
rect 110644 176972 110708 176976
rect 123156 176972 123220 177036
rect 127020 176972 127084 177036
rect 101996 176836 102060 176900
rect 104572 176760 104636 176764
rect 104572 176704 104622 176760
rect 104622 176704 104636 176760
rect 104572 176700 104636 176704
rect 108068 176760 108132 176764
rect 108068 176704 108118 176760
rect 108118 176704 108132 176760
rect 108068 176700 108132 176704
rect 109540 176700 109604 176764
rect 115796 176760 115860 176764
rect 115796 176704 115846 176760
rect 115846 176704 115860 176760
rect 115796 176700 115860 176704
rect 124444 176760 124508 176764
rect 124444 176704 124494 176760
rect 124494 176704 124508 176760
rect 124444 176700 124508 176704
rect 125732 176700 125796 176764
rect 130700 176760 130764 176764
rect 130700 176704 130750 176760
rect 130750 176704 130764 176760
rect 130700 176700 130764 176704
rect 134380 176700 134444 176764
rect 136036 176760 136100 176764
rect 136036 176704 136086 176760
rect 136086 176704 136100 176760
rect 136036 176700 136100 176704
rect 148180 176760 148244 176764
rect 148180 176704 148230 176760
rect 148230 176704 148244 176760
rect 148180 176700 148244 176704
rect 260052 176700 260116 176764
rect 99420 176428 99484 176492
rect 103284 176428 103348 176492
rect 249196 176020 249260 176084
rect 260972 175884 261036 175948
rect 100708 175400 100772 175404
rect 100708 175344 100758 175400
rect 100758 175344 100772 175400
rect 100708 175340 100772 175344
rect 121868 175400 121932 175404
rect 121868 175344 121918 175400
rect 121918 175344 121932 175400
rect 121868 175340 121932 175344
rect 128124 175400 128188 175404
rect 128124 175344 128174 175400
rect 128174 175344 128188 175400
rect 128124 175340 128188 175344
rect 158852 175400 158916 175404
rect 158852 175344 158902 175400
rect 158902 175344 158916 175400
rect 158852 175340 158916 175344
rect 262812 175340 262876 175404
rect 113142 174992 113206 174996
rect 113142 174936 113178 174992
rect 113178 174936 113206 174992
rect 113142 174932 113206 174936
rect 119398 174992 119462 174996
rect 119398 174936 119434 174992
rect 119434 174936 119462 174992
rect 119398 174932 119462 174936
rect 249196 174252 249260 174316
rect 249380 173300 249444 173364
rect 321324 170580 321388 170644
rect 260972 170308 261036 170372
rect 338620 165684 338684 165748
rect 254532 163372 254596 163436
rect 166396 161468 166460 161532
rect 259500 160788 259564 160852
rect 269068 157388 269132 157452
rect 258396 155212 258460 155276
rect 166212 154532 166276 154596
rect 258580 153444 258644 153508
rect 266308 153308 266372 153372
rect 251772 148140 251836 148204
rect 255268 147460 255332 147524
rect 307708 146372 307772 146436
rect 258396 146236 258460 146300
rect 307708 145556 307772 145620
rect 263548 144468 263612 144532
rect 168972 142156 169036 142220
rect 251956 142292 252020 142356
rect 267780 140796 267844 140860
rect 256740 140388 256804 140452
rect 263732 138756 263796 138820
rect 342116 138076 342180 138140
rect 166212 135492 166276 135556
rect 336780 135220 336844 135284
rect 302740 133996 302804 134060
rect 251956 130868 252020 130932
rect 305500 130052 305564 130116
rect 170260 128556 170324 128620
rect 173020 127196 173084 127260
rect 169156 127060 169220 127124
rect 299980 118084 300044 118148
rect 166948 115832 167012 115836
rect 166948 115776 166962 115832
rect 166962 115776 167012 115832
rect 166948 115772 167012 115776
rect 335492 115908 335556 115972
rect 331444 114684 331508 114748
rect 345060 114548 345124 114612
rect 307156 114004 307220 114068
rect 301820 113460 301884 113524
rect 258580 112916 258644 112980
rect 251772 112644 251836 112708
rect 302924 112100 302988 112164
rect 332548 110604 332612 110668
rect 338252 110468 338316 110532
rect 334204 109516 334268 109580
rect 335124 109108 335188 109172
rect 327212 107748 327276 107812
rect 342300 106388 342364 106452
rect 327028 106252 327092 106316
rect 214420 105164 214484 105228
rect 304212 104076 304276 104140
rect 170444 102172 170508 102236
rect 304396 101900 304460 101964
rect 334020 100948 334084 101012
rect 324268 100812 324332 100876
rect 305684 99588 305748 99652
rect 340092 99452 340156 99516
rect 166948 98016 167012 98020
rect 331260 98092 331324 98156
rect 166948 97960 166962 98016
rect 166962 97960 167012 98016
rect 166948 97956 167012 97960
rect 298692 97684 298756 97748
rect 166396 97140 166460 97204
rect 306972 97004 307036 97068
rect 262812 96732 262876 96796
rect 260052 96596 260116 96660
rect 166948 95100 167012 95164
rect 111918 94692 111982 94756
rect 113686 94752 113750 94756
rect 113686 94696 113730 94752
rect 113730 94696 113750 94752
rect 113686 94692 113750 94696
rect 129326 94752 129390 94756
rect 129326 94696 129370 94752
rect 129370 94696 129390 94752
rect 129326 94692 129390 94696
rect 151630 94752 151694 94756
rect 151630 94696 151634 94752
rect 151634 94696 151690 94752
rect 151690 94696 151694 94752
rect 151630 94692 151694 94696
rect 214420 93740 214484 93804
rect 118004 93664 118068 93668
rect 118004 93608 118054 93664
rect 118054 93608 118068 93664
rect 118004 93604 118068 93608
rect 133092 93664 133156 93668
rect 133092 93608 133142 93664
rect 133142 93608 133156 93664
rect 133092 93604 133156 93608
rect 85620 93528 85684 93532
rect 85620 93472 85670 93528
rect 85670 93472 85684 93528
rect 85620 93468 85684 93472
rect 107700 93528 107764 93532
rect 107700 93472 107750 93528
rect 107750 93472 107764 93528
rect 107700 93468 107764 93472
rect 120580 93528 120644 93532
rect 120580 93472 120630 93528
rect 120630 93472 120644 93528
rect 120580 93468 120644 93472
rect 110092 93256 110156 93260
rect 110092 93200 110142 93256
rect 110142 93200 110156 93256
rect 110092 93196 110156 93200
rect 84332 92380 84396 92444
rect 91324 92380 91388 92444
rect 95004 92440 95068 92444
rect 95004 92384 95054 92440
rect 95054 92384 95068 92440
rect 95004 92380 95068 92384
rect 105676 92380 105740 92444
rect 115428 92440 115492 92444
rect 115428 92384 115478 92440
rect 115478 92384 115492 92440
rect 115428 92380 115492 92384
rect 116716 92440 116780 92444
rect 116716 92384 116766 92440
rect 116766 92384 116780 92440
rect 116716 92380 116780 92384
rect 120212 92380 120276 92444
rect 125364 92380 125428 92444
rect 125916 92440 125980 92444
rect 125916 92384 125966 92440
rect 125966 92384 125980 92440
rect 125916 92380 125980 92384
rect 130700 92440 130764 92444
rect 130700 92384 130750 92440
rect 130750 92384 130764 92440
rect 130700 92380 130764 92384
rect 151676 92440 151740 92444
rect 151676 92384 151726 92440
rect 151726 92384 151740 92440
rect 151676 92380 151740 92384
rect 152044 92440 152108 92444
rect 152044 92384 152094 92440
rect 152094 92384 152108 92440
rect 152044 92380 152108 92384
rect 109172 92244 109236 92308
rect 119292 92244 119356 92308
rect 166396 92244 166460 92308
rect 136036 92108 136100 92172
rect 90220 91700 90284 91764
rect 102548 91700 102612 91764
rect 114876 91700 114940 91764
rect 126652 91760 126716 91764
rect 126652 91704 126702 91760
rect 126702 91704 126716 91760
rect 126652 91700 126716 91704
rect 99972 91624 100036 91628
rect 99972 91568 100022 91624
rect 100022 91568 100036 91624
rect 99972 91564 100036 91568
rect 102732 91564 102796 91628
rect 98132 91428 98196 91492
rect 101812 91488 101876 91492
rect 101812 91432 101862 91488
rect 101862 91432 101876 91488
rect 101812 91428 101876 91432
rect 122788 91488 122852 91492
rect 122788 91432 122838 91488
rect 122838 91432 122852 91488
rect 122788 91428 122852 91432
rect 151124 91428 151188 91492
rect 96660 91292 96724 91356
rect 98500 91292 98564 91356
rect 100892 91292 100956 91356
rect 106412 91292 106476 91356
rect 111196 91292 111260 91356
rect 114324 91352 114388 91356
rect 114324 91296 114374 91352
rect 114374 91296 114388 91352
rect 114324 91292 114388 91296
rect 121684 91292 121748 91356
rect 74764 91156 74828 91220
rect 86724 91156 86788 91220
rect 88012 91216 88076 91220
rect 88012 91160 88062 91216
rect 88062 91160 88076 91216
rect 88012 91156 88076 91160
rect 88932 91156 88996 91220
rect 92612 91156 92676 91220
rect 93900 91156 93964 91220
rect 96292 91156 96356 91220
rect 97212 91156 97276 91220
rect 99052 91156 99116 91220
rect 100524 91216 100588 91220
rect 100524 91160 100574 91216
rect 100574 91160 100588 91216
rect 100524 91156 100588 91160
rect 101996 91216 102060 91220
rect 101996 91160 102010 91216
rect 102010 91160 102060 91216
rect 101996 91156 102060 91160
rect 104204 91216 104268 91220
rect 104204 91160 104254 91216
rect 104254 91160 104268 91216
rect 104204 91156 104268 91160
rect 104572 91156 104636 91220
rect 105492 91156 105556 91220
rect 106780 91156 106844 91220
rect 108068 91156 108132 91220
rect 109540 91216 109604 91220
rect 109540 91160 109590 91216
rect 109590 91160 109604 91216
rect 109540 91156 109604 91160
rect 110644 91156 110708 91220
rect 112300 91216 112364 91220
rect 112300 91160 112350 91216
rect 112350 91160 112364 91216
rect 112300 91156 112364 91160
rect 113220 91156 113284 91220
rect 115796 91216 115860 91220
rect 115796 91160 115846 91216
rect 115846 91160 115860 91216
rect 115796 91156 115860 91160
rect 117084 91216 117148 91220
rect 117084 91160 117134 91216
rect 117134 91160 117148 91216
rect 117084 91156 117148 91160
rect 118188 91156 118252 91220
rect 119660 91156 119724 91220
rect 122052 91156 122116 91220
rect 123156 91156 123220 91220
rect 124076 91216 124140 91220
rect 124076 91160 124126 91216
rect 124126 91160 124140 91216
rect 124076 91156 124140 91160
rect 124444 91156 124508 91220
rect 126468 91216 126532 91220
rect 126468 91160 126518 91216
rect 126518 91160 126532 91216
rect 126468 91156 126532 91160
rect 127572 91156 127636 91220
rect 132356 91216 132420 91220
rect 132356 91160 132406 91216
rect 132406 91160 132420 91216
rect 132356 91156 132420 91160
rect 134380 91156 134444 91220
rect 170444 91020 170508 91084
rect 168972 89660 169036 89724
rect 166212 88164 166276 88228
rect 173020 81364 173084 81428
rect 170260 80004 170324 80068
rect 169156 78508 169220 78572
rect 304396 62732 304460 62796
rect 302924 61372 302988 61436
rect 298692 57156 298756 57220
rect 301820 54436 301884 54500
rect 305500 47500 305564 47564
rect 307156 32404 307220 32468
rect 299980 30908 300044 30972
rect 302740 29548 302804 29612
rect 305684 18532 305748 18596
rect 304212 12956 304276 13020
rect 306972 4796 307036 4860
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 59123 700364 59189 700365
rect 59123 700300 59124 700364
rect 59188 700300 59189 700364
rect 59123 700299 59189 700300
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 59126 241773 59186 700299
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 61883 456924 61949 456925
rect 61883 456860 61884 456924
rect 61948 456860 61949 456924
rect 61883 456859 61949 456860
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59123 241772 59189 241773
rect 59123 241708 59124 241772
rect 59188 241708 59189 241772
rect 59123 241707 59189 241708
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 61886 240413 61946 456859
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 70899 702540 70965 702541
rect 70899 702476 70900 702540
rect 70964 702476 70965 702540
rect 70899 702475 70965 702476
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 68875 313988 68941 313989
rect 68875 313924 68876 313988
rect 68940 313924 68941 313988
rect 68875 313923 68941 313924
rect 68878 288421 68938 313923
rect 70902 296730 70962 702475
rect 70534 296670 70962 296730
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 70534 288829 70594 296670
rect 73794 294000 74414 326898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 294000 78134 294618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 294000 81854 298338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 294000 85574 302058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 294000 92414 308898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 385174 96134 420618
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 313174 96134 348618
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 294000 96134 312618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 424894 99854 460338
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 388894 99854 424338
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 352894 99854 388338
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 294000 99854 316338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 356614 103574 392058
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 320614 103574 356058
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 294000 103574 320058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 294000 110414 326898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 294000 114134 294618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 294000 117854 298338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 294000 121574 302058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 120027 293996 120093 293997
rect 120027 293932 120028 293996
rect 120092 293932 120093 293996
rect 120027 293931 120093 293932
rect 120030 289237 120090 293931
rect 120027 289236 120093 289237
rect 120027 289172 120028 289236
rect 120092 289172 120093 289236
rect 120027 289171 120093 289172
rect 70531 288828 70597 288829
rect 70531 288764 70532 288828
rect 70596 288764 70597 288828
rect 70531 288763 70597 288764
rect 68875 288420 68941 288421
rect 68875 288356 68876 288420
rect 68940 288356 68941 288420
rect 68875 288355 68941 288356
rect 122051 287740 122117 287741
rect 122051 287676 122052 287740
rect 122116 287676 122117 287740
rect 122051 287675 122117 287676
rect 64643 284476 64709 284477
rect 64643 284412 64644 284476
rect 64708 284412 64709 284476
rect 64643 284411 64709 284412
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 62987 254148 63053 254149
rect 62987 254084 62988 254148
rect 63052 254084 63053 254148
rect 62987 254083 63053 254084
rect 61883 240412 61949 240413
rect 61883 240348 61884 240412
rect 61948 240348 61949 240412
rect 61883 240347 61949 240348
rect 62990 232525 63050 254083
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 62987 232524 63053 232525
rect 62987 232460 62988 232524
rect 63052 232460 63053 232524
rect 62987 232459 63053 232460
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 208894 63854 244338
rect 64646 226949 64706 284411
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66115 256732 66181 256733
rect 66115 256668 66116 256732
rect 66180 256668 66181 256732
rect 66115 256667 66181 256668
rect 66118 236605 66178 256667
rect 66954 248614 67574 284058
rect 89568 273454 89888 273486
rect 89568 273218 89610 273454
rect 89846 273218 89888 273454
rect 89568 273134 89888 273218
rect 89568 272898 89610 273134
rect 89846 272898 89888 273134
rect 89568 272866 89888 272898
rect 122054 269789 122114 287675
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 122051 269788 122117 269789
rect 122051 269724 122052 269788
rect 122116 269724 122117 269788
rect 122051 269723 122117 269724
rect 74208 255454 74528 255486
rect 74208 255218 74250 255454
rect 74486 255218 74528 255454
rect 74208 255134 74528 255218
rect 74208 254898 74250 255134
rect 74486 254898 74528 255134
rect 74208 254866 74528 254898
rect 104928 255454 105248 255486
rect 104928 255218 104970 255454
rect 105206 255218 105248 255454
rect 104928 255134 105248 255218
rect 104928 254898 104970 255134
rect 105206 254898 105248 255134
rect 104928 254866 105248 254898
rect 120027 253196 120093 253197
rect 120027 253132 120028 253196
rect 120092 253132 120093 253196
rect 120027 253131 120093 253132
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66115 236604 66181 236605
rect 66115 236540 66116 236604
rect 66180 236540 66181 236604
rect 66115 236539 66181 236540
rect 64643 226948 64709 226949
rect 64643 226884 64644 226948
rect 64708 226884 64709 226948
rect 64643 226883 64709 226884
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 66954 212614 67574 248058
rect 120030 239869 120090 253131
rect 120027 239868 120093 239869
rect 120027 239804 120028 239868
rect 120092 239804 120093 239868
rect 120027 239803 120093 239804
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176600 67574 212058
rect 73794 219454 74414 238000
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 176600 74414 182898
rect 77514 223174 78134 238000
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 176600 78134 186618
rect 81234 226894 81854 238000
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 176600 81854 190338
rect 84954 230614 85574 238000
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 176600 85574 194058
rect 91794 237454 92414 238000
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 176600 92414 200898
rect 95514 205174 96134 238000
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 176600 96134 204618
rect 99234 208894 99854 238000
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 97027 177716 97093 177717
rect 97027 177652 97028 177716
rect 97092 177652 97093 177716
rect 97027 177651 97093 177652
rect 98315 177716 98381 177717
rect 98315 177652 98316 177716
rect 98380 177652 98381 177716
rect 98315 177651 98381 177652
rect 97030 175130 97090 177651
rect 96960 175070 97090 175130
rect 98318 175130 98378 177651
rect 99234 176600 99854 208338
rect 102954 212614 103574 238000
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 101995 176900 102061 176901
rect 101995 176836 101996 176900
rect 102060 176836 102061 176900
rect 101995 176835 102061 176836
rect 99419 176492 99485 176493
rect 99419 176428 99420 176492
rect 99484 176428 99485 176492
rect 99419 176427 99485 176428
rect 99422 175130 99482 176427
rect 100707 175404 100773 175405
rect 100707 175340 100708 175404
rect 100772 175340 100773 175404
rect 100707 175339 100773 175340
rect 98318 175070 98380 175130
rect 96960 174494 97020 175070
rect 98320 174494 98380 175070
rect 99408 175070 99482 175130
rect 100710 175130 100770 175339
rect 101998 175130 102058 176835
rect 102954 176600 103574 212058
rect 109794 219454 110414 238000
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 105675 177716 105741 177717
rect 105675 177652 105676 177716
rect 105740 177652 105741 177716
rect 105675 177651 105741 177652
rect 106963 177716 107029 177717
rect 106963 177652 106964 177716
rect 107028 177652 107029 177716
rect 106963 177651 107029 177652
rect 104571 176764 104637 176765
rect 104571 176700 104572 176764
rect 104636 176700 104637 176764
rect 104571 176699 104637 176700
rect 103283 176492 103349 176493
rect 103283 176428 103284 176492
rect 103348 176428 103349 176492
rect 103283 176427 103349 176428
rect 100710 175070 100828 175130
rect 99408 174494 99468 175070
rect 100768 174494 100828 175070
rect 101992 175070 102058 175130
rect 103286 175130 103346 176427
rect 104574 175130 104634 176699
rect 105678 175130 105738 177651
rect 103286 175070 103412 175130
rect 104574 175070 104636 175130
rect 101992 174494 102052 175070
rect 103352 174494 103412 175070
rect 104576 174494 104636 175070
rect 105664 175070 105738 175130
rect 106966 175130 107026 177651
rect 108067 176764 108133 176765
rect 108067 176700 108068 176764
rect 108132 176700 108133 176764
rect 108067 176699 108133 176700
rect 109539 176764 109605 176765
rect 109539 176700 109540 176764
rect 109604 176700 109605 176764
rect 109539 176699 109605 176700
rect 108070 175130 108130 176699
rect 106966 175070 107084 175130
rect 108070 175070 108172 175130
rect 105664 174494 105724 175070
rect 107024 174494 107084 175070
rect 108112 174494 108172 175070
rect 109542 174994 109602 176699
rect 109794 176600 110414 182898
rect 113514 223174 114134 238000
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 112115 177172 112181 177173
rect 112115 177108 112116 177172
rect 112180 177108 112181 177172
rect 112115 177107 112181 177108
rect 110643 177036 110709 177037
rect 110643 176972 110644 177036
rect 110708 176972 110709 177036
rect 110643 176971 110709 176972
rect 110646 175130 110706 176971
rect 112118 175130 112178 177107
rect 113514 176600 114134 186618
rect 117234 226894 117854 238000
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 114323 177716 114389 177717
rect 114323 177652 114324 177716
rect 114388 177652 114389 177716
rect 114323 177651 114389 177652
rect 116899 177716 116965 177717
rect 116899 177652 116900 177716
rect 116964 177652 116965 177716
rect 116899 177651 116965 177652
rect 110646 175070 110756 175130
rect 109472 174934 109602 174994
rect 109472 174494 109532 174934
rect 110696 174494 110756 175070
rect 112056 175070 112178 175130
rect 114326 175130 114386 177651
rect 115795 176764 115861 176765
rect 115795 176700 115796 176764
rect 115860 176700 115861 176764
rect 115795 176699 115861 176700
rect 115798 175130 115858 176699
rect 114326 175070 114428 175130
rect 112056 174494 112116 175070
rect 113141 174996 113207 174997
rect 113141 174932 113142 174996
rect 113206 174932 113207 174996
rect 113141 174931 113207 174932
rect 113144 174494 113204 174931
rect 114368 174494 114428 175070
rect 115728 175070 115858 175130
rect 116902 175130 116962 177651
rect 117234 176600 117854 190338
rect 120954 230614 121574 238000
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 118371 177716 118437 177717
rect 118371 177652 118372 177716
rect 118436 177652 118437 177716
rect 118371 177651 118437 177652
rect 120763 177716 120829 177717
rect 120763 177652 120764 177716
rect 120828 177652 120829 177716
rect 120763 177651 120829 177652
rect 118374 175130 118434 177651
rect 120766 175130 120826 177651
rect 120954 176600 121574 194058
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 123155 177036 123221 177037
rect 123155 176972 123156 177036
rect 123220 176972 123221 177036
rect 123155 176971 123221 176972
rect 127019 177036 127085 177037
rect 127019 176972 127020 177036
rect 127084 176972 127085 177036
rect 127019 176971 127085 176972
rect 121867 175404 121933 175405
rect 121867 175340 121868 175404
rect 121932 175340 121933 175404
rect 121867 175339 121933 175340
rect 121870 175130 121930 175339
rect 123158 175130 123218 176971
rect 124443 176764 124509 176765
rect 124443 176700 124444 176764
rect 124508 176700 124509 176764
rect 124443 176699 124509 176700
rect 125731 176764 125797 176765
rect 125731 176700 125732 176764
rect 125796 176700 125797 176764
rect 125731 176699 125797 176700
rect 124446 175130 124506 176699
rect 125734 175130 125794 176699
rect 127022 175130 127082 176971
rect 127794 176600 128414 200898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 129411 177716 129477 177717
rect 129411 177652 129412 177716
rect 129476 177652 129477 177716
rect 129411 177651 129477 177652
rect 128123 175404 128189 175405
rect 128123 175340 128124 175404
rect 128188 175340 128189 175404
rect 128123 175339 128189 175340
rect 128126 175130 128186 175339
rect 116902 175070 117012 175130
rect 115728 174494 115788 175070
rect 116952 174494 117012 175070
rect 118312 175070 118434 175130
rect 120760 175070 120826 175130
rect 121848 175070 121930 175130
rect 123072 175070 123218 175130
rect 124432 175070 124506 175130
rect 125656 175070 125794 175130
rect 127016 175070 127082 175130
rect 128104 175070 128186 175130
rect 129414 175130 129474 177651
rect 130699 176764 130765 176765
rect 130699 176700 130700 176764
rect 130764 176700 130765 176764
rect 130699 176699 130765 176700
rect 130702 175130 130762 176699
rect 131514 176600 132134 204618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 132355 177716 132421 177717
rect 132355 177652 132356 177716
rect 132420 177652 132421 177716
rect 132355 177651 132421 177652
rect 133091 177716 133157 177717
rect 133091 177652 133092 177716
rect 133156 177652 133157 177716
rect 133091 177651 133157 177652
rect 132358 175130 132418 177651
rect 129414 175070 129524 175130
rect 118312 174494 118372 175070
rect 119397 174996 119463 174997
rect 119397 174932 119398 174996
rect 119462 174932 119463 174996
rect 119397 174931 119463 174932
rect 119400 174494 119460 174931
rect 120760 174494 120820 175070
rect 121848 174494 121908 175070
rect 123072 174494 123132 175070
rect 124432 174494 124492 175070
rect 125656 174494 125716 175070
rect 127016 174494 127076 175070
rect 128104 174494 128164 175070
rect 129464 174494 129524 175070
rect 130688 175070 130762 175130
rect 132048 175070 132418 175130
rect 133094 175130 133154 177651
rect 134379 176764 134445 176765
rect 134379 176700 134380 176764
rect 134444 176700 134445 176764
rect 134379 176699 134445 176700
rect 134382 175130 134442 176699
rect 135234 176600 135854 208338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 136035 176764 136101 176765
rect 136035 176700 136036 176764
rect 136100 176700 136101 176764
rect 136035 176699 136101 176700
rect 136038 175130 136098 176699
rect 138954 176600 139574 212058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 176600 146414 182898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 148179 176764 148245 176765
rect 148179 176700 148180 176764
rect 148244 176700 148245 176764
rect 148179 176699 148245 176700
rect 133094 175070 133196 175130
rect 130688 174494 130748 175070
rect 132048 174494 132108 175070
rect 133136 174494 133196 175070
rect 134360 175070 134442 175130
rect 135720 175070 136098 175130
rect 148182 175130 148242 176699
rect 149514 176600 150134 186618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 176600 153854 190338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 176600 157574 194058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 166947 271964 167013 271965
rect 166947 271900 166948 271964
rect 167012 271900 167013 271964
rect 166947 271899 167013 271900
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 176600 164414 200898
rect 166211 183700 166277 183701
rect 166211 183636 166212 183700
rect 166276 183636 166277 183700
rect 166211 183635 166277 183636
rect 158851 175404 158917 175405
rect 158851 175340 158852 175404
rect 158916 175340 158917 175404
rect 158851 175339 158917 175340
rect 158854 175130 158914 175339
rect 148182 175070 148292 175130
rect 134360 174494 134420 175070
rect 135720 174494 135780 175070
rect 148232 174494 148292 175070
rect 158840 175070 158914 175130
rect 158840 174494 158900 175070
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 69072 165454 69420 165486
rect 69072 165218 69128 165454
rect 69364 165218 69420 165454
rect 69072 165134 69420 165218
rect 69072 164898 69128 165134
rect 69364 164898 69420 165134
rect 69072 164866 69420 164898
rect 164136 165454 164484 165486
rect 164136 165218 164192 165454
rect 164428 165218 164484 165454
rect 164136 165134 164484 165218
rect 164136 164898 164192 165134
rect 164428 164898 164484 165134
rect 164136 164866 164484 164898
rect 166214 154597 166274 183635
rect 166395 179484 166461 179485
rect 166395 179420 166396 179484
rect 166460 179420 166461 179484
rect 166395 179419 166461 179420
rect 166398 161533 166458 179419
rect 166395 161532 166461 161533
rect 166395 161468 166396 161532
rect 166460 161468 166461 161532
rect 166395 161467 166461 161468
rect 166211 154596 166277 154597
rect 166211 154532 166212 154596
rect 166276 154532 166277 154596
rect 166211 154531 166277 154532
rect 69752 147454 70100 147486
rect 69752 147218 69808 147454
rect 70044 147218 70100 147454
rect 69752 147134 70100 147218
rect 69752 146898 69808 147134
rect 70044 146898 70100 147134
rect 69752 146866 70100 146898
rect 163456 147454 163804 147486
rect 163456 147218 163512 147454
rect 163748 147218 163804 147454
rect 163456 147134 163804 147218
rect 163456 146898 163512 147134
rect 163748 146898 163804 147134
rect 163456 146866 163804 146898
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 166211 135556 166277 135557
rect 166211 135492 166212 135556
rect 166276 135492 166277 135556
rect 166211 135491 166277 135492
rect 69072 129454 69420 129486
rect 69072 129218 69128 129454
rect 69364 129218 69420 129454
rect 69072 129134 69420 129218
rect 69072 128898 69128 129134
rect 69364 128898 69420 129134
rect 69072 128866 69420 128898
rect 164136 129454 164484 129486
rect 164136 129218 164192 129454
rect 164428 129218 164484 129454
rect 164136 129134 164484 129218
rect 164136 128898 164192 129134
rect 164428 128898 164484 129134
rect 164136 128866 164484 128898
rect 69752 111454 70100 111486
rect 69752 111218 69808 111454
rect 70044 111218 70100 111454
rect 69752 111134 70100 111218
rect 69752 110898 69808 111134
rect 70044 110898 70100 111134
rect 69752 110866 70100 110898
rect 163456 111454 163804 111486
rect 163456 111218 163512 111454
rect 163748 111218 163804 111454
rect 163456 111134 163804 111218
rect 163456 110898 163512 111134
rect 163748 110898 163804 111134
rect 163456 110866 163804 110898
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 74656 94890 74716 95200
rect 84312 94890 84372 95200
rect 85536 94890 85596 95200
rect 86624 94890 86684 95200
rect 87984 94890 88044 95200
rect 88936 94890 88996 95200
rect 74656 94830 74826 94890
rect 84312 94830 84394 94890
rect 85536 94830 85682 94890
rect 86624 94830 86786 94890
rect 87984 94830 88074 94890
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 68614 67574 93100
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 75454 74414 93100
rect 74766 91221 74826 94830
rect 74763 91220 74829 91221
rect 74763 91156 74764 91220
rect 74828 91156 74829 91220
rect 74763 91155 74829 91156
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 79174 78134 93100
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 82894 81854 93100
rect 84334 92445 84394 94830
rect 85622 93533 85682 94830
rect 85619 93532 85685 93533
rect 85619 93468 85620 93532
rect 85684 93468 85685 93532
rect 85619 93467 85685 93468
rect 84331 92444 84397 92445
rect 84331 92380 84332 92444
rect 84396 92380 84397 92444
rect 84331 92379 84397 92380
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 86614 85574 93100
rect 86726 91221 86786 94830
rect 88014 91221 88074 94830
rect 88934 94830 88996 94890
rect 90160 94890 90220 95200
rect 91384 94890 91444 95200
rect 90160 94830 90282 94890
rect 88934 91221 88994 94830
rect 90222 91765 90282 94830
rect 91326 94830 91444 94890
rect 92472 94890 92532 95200
rect 93832 94890 93892 95200
rect 94920 94890 94980 95200
rect 96008 94890 96068 95200
rect 96688 94890 96748 95200
rect 92472 94830 92674 94890
rect 93832 94830 93962 94890
rect 94920 94830 95066 94890
rect 96008 94830 96354 94890
rect 91326 92445 91386 94830
rect 91323 92444 91389 92445
rect 91323 92380 91324 92444
rect 91388 92380 91389 92444
rect 91323 92379 91389 92380
rect 90219 91764 90285 91765
rect 90219 91700 90220 91764
rect 90284 91700 90285 91764
rect 90219 91699 90285 91700
rect 86723 91220 86789 91221
rect 86723 91156 86724 91220
rect 86788 91156 86789 91220
rect 86723 91155 86789 91156
rect 88011 91220 88077 91221
rect 88011 91156 88012 91220
rect 88076 91156 88077 91220
rect 88011 91155 88077 91156
rect 88931 91220 88997 91221
rect 88931 91156 88932 91220
rect 88996 91156 88997 91220
rect 88931 91155 88997 91156
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 93100
rect 92614 91221 92674 94830
rect 93902 91221 93962 94830
rect 95006 92445 95066 94830
rect 95003 92444 95069 92445
rect 95003 92380 95004 92444
rect 95068 92380 95069 92444
rect 95003 92379 95069 92380
rect 92611 91220 92677 91221
rect 92611 91156 92612 91220
rect 92676 91156 92677 91220
rect 92611 91155 92677 91156
rect 93899 91220 93965 91221
rect 93899 91156 93900 91220
rect 93964 91156 93965 91220
rect 93899 91155 93965 91156
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 61174 96134 93100
rect 96294 91221 96354 94830
rect 96662 94830 96748 94890
rect 97096 94890 97156 95200
rect 98048 94890 98108 95200
rect 98456 94890 98516 95200
rect 99136 94890 99196 95200
rect 97096 94830 97274 94890
rect 98048 94830 98194 94890
rect 98456 94830 98562 94890
rect 96662 91357 96722 94830
rect 96659 91356 96725 91357
rect 96659 91292 96660 91356
rect 96724 91292 96725 91356
rect 96659 91291 96725 91292
rect 97214 91221 97274 94830
rect 98134 91493 98194 94830
rect 98131 91492 98197 91493
rect 98131 91428 98132 91492
rect 98196 91428 98197 91492
rect 98131 91427 98197 91428
rect 98502 91357 98562 94830
rect 99054 94830 99196 94890
rect 99544 94890 99604 95200
rect 100632 94890 100692 95200
rect 99544 94830 100034 94890
rect 98499 91356 98565 91357
rect 98499 91292 98500 91356
rect 98564 91292 98565 91356
rect 98499 91291 98565 91292
rect 99054 91221 99114 94830
rect 96291 91220 96357 91221
rect 96291 91156 96292 91220
rect 96356 91156 96357 91220
rect 96291 91155 96357 91156
rect 97211 91220 97277 91221
rect 97211 91156 97212 91220
rect 97276 91156 97277 91220
rect 97211 91155 97277 91156
rect 99051 91220 99117 91221
rect 99051 91156 99052 91220
rect 99116 91156 99117 91220
rect 99051 91155 99117 91156
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 64894 99854 93100
rect 99974 91629 100034 94830
rect 100526 94830 100692 94890
rect 100768 94890 100828 95200
rect 101856 94890 101916 95200
rect 100768 94830 100954 94890
rect 99971 91628 100037 91629
rect 99971 91564 99972 91628
rect 100036 91564 100037 91628
rect 99971 91563 100037 91564
rect 100526 91221 100586 94830
rect 100894 91357 100954 94830
rect 101814 94830 101916 94890
rect 101992 94890 102052 95200
rect 102944 94890 103004 95200
rect 103216 94890 103276 95200
rect 104304 94890 104364 95200
rect 101992 94830 102058 94890
rect 101814 91493 101874 94830
rect 101811 91492 101877 91493
rect 101811 91428 101812 91492
rect 101876 91428 101877 91492
rect 101811 91427 101877 91428
rect 100891 91356 100957 91357
rect 100891 91292 100892 91356
rect 100956 91292 100957 91356
rect 100891 91291 100957 91292
rect 101998 91221 102058 94830
rect 102550 94830 103004 94890
rect 103102 94830 103276 94890
rect 104206 94830 104364 94890
rect 104440 94890 104500 95200
rect 105392 94890 105452 95200
rect 105664 94890 105724 95200
rect 106480 94890 106540 95200
rect 104440 94830 104634 94890
rect 105392 94830 105554 94890
rect 105664 94830 105738 94890
rect 102550 91765 102610 94830
rect 103102 93870 103162 94830
rect 102734 93810 103162 93870
rect 102547 91764 102613 91765
rect 102547 91700 102548 91764
rect 102612 91700 102613 91764
rect 102547 91699 102613 91700
rect 102734 91629 102794 93810
rect 102731 91628 102797 91629
rect 102731 91564 102732 91628
rect 102796 91564 102797 91628
rect 102731 91563 102797 91564
rect 100523 91220 100589 91221
rect 100523 91156 100524 91220
rect 100588 91156 100589 91220
rect 100523 91155 100589 91156
rect 101995 91220 102061 91221
rect 101995 91156 101996 91220
rect 102060 91156 102061 91220
rect 101995 91155 102061 91156
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 68614 103574 93100
rect 104206 91221 104266 94830
rect 104574 91221 104634 94830
rect 105494 91221 105554 94830
rect 105678 92445 105738 94830
rect 106414 94830 106540 94890
rect 106616 94890 106676 95200
rect 107704 94890 107764 95200
rect 108112 94890 108172 95200
rect 106616 94830 106842 94890
rect 105675 92444 105741 92445
rect 105675 92380 105676 92444
rect 105740 92380 105741 92444
rect 105675 92379 105741 92380
rect 106414 91357 106474 94830
rect 106411 91356 106477 91357
rect 106411 91292 106412 91356
rect 106476 91292 106477 91356
rect 106411 91291 106477 91292
rect 106782 91221 106842 94830
rect 107702 94830 107764 94890
rect 108070 94830 108172 94890
rect 109064 94890 109124 95200
rect 109472 94890 109532 95200
rect 110152 94890 110212 95200
rect 110696 94890 110756 95200
rect 111240 94890 111300 95200
rect 109064 94830 109234 94890
rect 109472 94830 109602 94890
rect 107702 93533 107762 94830
rect 107699 93532 107765 93533
rect 107699 93468 107700 93532
rect 107764 93468 107765 93532
rect 107699 93467 107765 93468
rect 108070 91221 108130 94830
rect 109174 92309 109234 94830
rect 109171 92308 109237 92309
rect 109171 92244 109172 92308
rect 109236 92244 109237 92308
rect 109171 92243 109237 92244
rect 109542 91221 109602 94830
rect 110094 94830 110212 94890
rect 110646 94830 110756 94890
rect 111198 94830 111300 94890
rect 110094 93261 110154 94830
rect 110091 93260 110157 93261
rect 110091 93196 110092 93260
rect 110156 93196 110157 93260
rect 110091 93195 110157 93196
rect 104203 91220 104269 91221
rect 104203 91156 104204 91220
rect 104268 91156 104269 91220
rect 104203 91155 104269 91156
rect 104571 91220 104637 91221
rect 104571 91156 104572 91220
rect 104636 91156 104637 91220
rect 104571 91155 104637 91156
rect 105491 91220 105557 91221
rect 105491 91156 105492 91220
rect 105556 91156 105557 91220
rect 105491 91155 105557 91156
rect 106779 91220 106845 91221
rect 106779 91156 106780 91220
rect 106844 91156 106845 91220
rect 106779 91155 106845 91156
rect 108067 91220 108133 91221
rect 108067 91156 108068 91220
rect 108132 91156 108133 91220
rect 108067 91155 108133 91156
rect 109539 91220 109605 91221
rect 109539 91156 109540 91220
rect 109604 91156 109605 91220
rect 109539 91155 109605 91156
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 75454 110414 93100
rect 110646 91221 110706 94830
rect 111198 91357 111258 94830
rect 111920 94757 111980 95200
rect 112328 94890 112388 95200
rect 112302 94830 112388 94890
rect 113144 94890 113204 95200
rect 113144 94830 113282 94890
rect 111917 94756 111983 94757
rect 111917 94692 111918 94756
rect 111982 94692 111983 94756
rect 111917 94691 111983 94692
rect 111195 91356 111261 91357
rect 111195 91292 111196 91356
rect 111260 91292 111261 91356
rect 111195 91291 111261 91292
rect 112302 91221 112362 94830
rect 113222 91221 113282 94830
rect 113688 94757 113748 95200
rect 114368 94890 114428 95200
rect 114326 94830 114428 94890
rect 114776 94890 114836 95200
rect 115456 94890 115516 95200
rect 115864 94890 115924 95200
rect 114776 94830 114938 94890
rect 113685 94756 113751 94757
rect 113685 94692 113686 94756
rect 113750 94692 113751 94756
rect 113685 94691 113751 94692
rect 110643 91220 110709 91221
rect 110643 91156 110644 91220
rect 110708 91156 110709 91220
rect 110643 91155 110709 91156
rect 112299 91220 112365 91221
rect 112299 91156 112300 91220
rect 112364 91156 112365 91220
rect 112299 91155 112365 91156
rect 113219 91220 113285 91221
rect 113219 91156 113220 91220
rect 113284 91156 113285 91220
rect 113219 91155 113285 91156
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 79174 114134 93100
rect 114326 91357 114386 94830
rect 114878 91765 114938 94830
rect 115430 94830 115516 94890
rect 115798 94830 115924 94890
rect 116680 94890 116740 95200
rect 117088 94890 117148 95200
rect 116680 94830 116778 94890
rect 115430 92445 115490 94830
rect 115427 92444 115493 92445
rect 115427 92380 115428 92444
rect 115492 92380 115493 92444
rect 115427 92379 115493 92380
rect 114875 91764 114941 91765
rect 114875 91700 114876 91764
rect 114940 91700 114941 91764
rect 114875 91699 114941 91700
rect 114323 91356 114389 91357
rect 114323 91292 114324 91356
rect 114388 91292 114389 91356
rect 114323 91291 114389 91292
rect 115798 91221 115858 94830
rect 116718 92445 116778 94830
rect 117086 94830 117148 94890
rect 117904 94890 117964 95200
rect 118176 94890 118236 95200
rect 119400 94890 119460 95200
rect 117904 94830 118066 94890
rect 118176 94830 118250 94890
rect 116715 92444 116781 92445
rect 116715 92380 116716 92444
rect 116780 92380 116781 92444
rect 116715 92379 116781 92380
rect 117086 91221 117146 94830
rect 118006 93669 118066 94830
rect 118003 93668 118069 93669
rect 118003 93604 118004 93668
rect 118068 93604 118069 93668
rect 118003 93603 118069 93604
rect 115795 91220 115861 91221
rect 115795 91156 115796 91220
rect 115860 91156 115861 91220
rect 115795 91155 115861 91156
rect 117083 91220 117149 91221
rect 117083 91156 117084 91220
rect 117148 91156 117149 91220
rect 117083 91155 117149 91156
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 82894 117854 93100
rect 118190 91221 118250 94830
rect 119294 94830 119460 94890
rect 119536 94890 119596 95200
rect 120216 94890 120276 95200
rect 120624 94890 120684 95200
rect 121712 94890 121772 95200
rect 119536 94830 119722 94890
rect 119294 92309 119354 94830
rect 119291 92308 119357 92309
rect 119291 92244 119292 92308
rect 119356 92244 119357 92308
rect 119291 92243 119357 92244
rect 119662 91221 119722 94830
rect 120214 94830 120276 94890
rect 120582 94830 120684 94890
rect 121686 94830 121772 94890
rect 121984 94890 122044 95200
rect 122800 94890 122860 95200
rect 123208 94890 123268 95200
rect 121984 94830 122114 94890
rect 122800 94830 123034 94890
rect 120214 92445 120274 94830
rect 120582 93533 120642 94830
rect 120579 93532 120645 93533
rect 120579 93468 120580 93532
rect 120644 93468 120645 93532
rect 120579 93467 120645 93468
rect 120211 92444 120277 92445
rect 120211 92380 120212 92444
rect 120276 92380 120277 92444
rect 120211 92379 120277 92380
rect 118187 91220 118253 91221
rect 118187 91156 118188 91220
rect 118252 91156 118253 91220
rect 118187 91155 118253 91156
rect 119659 91220 119725 91221
rect 119659 91156 119660 91220
rect 119724 91156 119725 91220
rect 119659 91155 119725 91156
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 86614 121574 93100
rect 121686 91357 121746 94830
rect 121683 91356 121749 91357
rect 121683 91292 121684 91356
rect 121748 91292 121749 91356
rect 121683 91291 121749 91292
rect 122054 91221 122114 94830
rect 122974 93870 123034 94830
rect 122606 93810 123034 93870
rect 123158 94830 123268 94890
rect 124024 94890 124084 95200
rect 124432 94890 124492 95200
rect 125384 94890 125444 95200
rect 124024 94830 124138 94890
rect 124432 94830 124506 94890
rect 122606 91490 122666 93810
rect 122787 91492 122853 91493
rect 122787 91490 122788 91492
rect 122606 91430 122788 91490
rect 122787 91428 122788 91430
rect 122852 91428 122853 91492
rect 122787 91427 122853 91428
rect 123158 91221 123218 94830
rect 124078 91221 124138 94830
rect 124446 91221 124506 94830
rect 125366 94830 125444 94890
rect 125656 94890 125716 95200
rect 126472 94890 126532 95200
rect 125656 94830 125978 94890
rect 125366 92445 125426 94830
rect 125918 92445 125978 94830
rect 126470 94830 126532 94890
rect 126608 94890 126668 95200
rect 128104 94890 128164 95200
rect 126608 94830 126714 94890
rect 125363 92444 125429 92445
rect 125363 92380 125364 92444
rect 125428 92380 125429 92444
rect 125363 92379 125429 92380
rect 125915 92444 125981 92445
rect 125915 92380 125916 92444
rect 125980 92380 125981 92444
rect 125915 92379 125981 92380
rect 126470 91221 126530 94830
rect 126654 91765 126714 94830
rect 127574 94830 128164 94890
rect 126651 91764 126717 91765
rect 126651 91700 126652 91764
rect 126716 91700 126717 91764
rect 126651 91699 126717 91700
rect 127574 91221 127634 94830
rect 129328 94757 129388 95200
rect 130688 94890 130748 95200
rect 131912 94890 131972 95200
rect 133136 94890 133196 95200
rect 130688 94830 130762 94890
rect 131912 94830 132418 94890
rect 129325 94756 129391 94757
rect 129325 94692 129326 94756
rect 129390 94692 129391 94756
rect 129325 94691 129391 94692
rect 122051 91220 122117 91221
rect 122051 91156 122052 91220
rect 122116 91156 122117 91220
rect 122051 91155 122117 91156
rect 123155 91220 123221 91221
rect 123155 91156 123156 91220
rect 123220 91156 123221 91220
rect 123155 91155 123221 91156
rect 124075 91220 124141 91221
rect 124075 91156 124076 91220
rect 124140 91156 124141 91220
rect 124075 91155 124141 91156
rect 124443 91220 124509 91221
rect 124443 91156 124444 91220
rect 124508 91156 124509 91220
rect 124443 91155 124509 91156
rect 126467 91220 126533 91221
rect 126467 91156 126468 91220
rect 126532 91156 126533 91220
rect 126467 91155 126533 91156
rect 127571 91220 127637 91221
rect 127571 91156 127572 91220
rect 127636 91156 127637 91220
rect 127571 91155 127637 91156
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 93100
rect 130702 92445 130762 94830
rect 130699 92444 130765 92445
rect 130699 92380 130700 92444
rect 130764 92380 130765 92444
rect 130699 92379 130765 92380
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 61174 132134 93100
rect 132358 91221 132418 94830
rect 133094 94830 133196 94890
rect 134360 94890 134420 95200
rect 135584 94890 135644 95200
rect 151496 94890 151556 95200
rect 134360 94830 134442 94890
rect 135584 94830 136098 94890
rect 133094 93669 133154 94830
rect 133091 93668 133157 93669
rect 133091 93604 133092 93668
rect 133156 93604 133157 93668
rect 133091 93603 133157 93604
rect 134382 91221 134442 94830
rect 132355 91220 132421 91221
rect 132355 91156 132356 91220
rect 132420 91156 132421 91220
rect 132355 91155 132421 91156
rect 134379 91220 134445 91221
rect 134379 91156 134380 91220
rect 134444 91156 134445 91220
rect 134379 91155 134445 91156
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 64894 135854 93100
rect 136038 92173 136098 94830
rect 151126 94830 151556 94890
rect 136035 92172 136101 92173
rect 136035 92108 136036 92172
rect 136100 92108 136101 92172
rect 136035 92107 136101 92108
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 68614 139574 93100
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 75454 146414 93100
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 79174 150134 93100
rect 151126 91493 151186 94830
rect 151632 94757 151692 95200
rect 151629 94756 151695 94757
rect 151629 94692 151630 94756
rect 151694 94692 151695 94756
rect 151629 94691 151695 94692
rect 151768 94210 151828 95200
rect 151904 94754 151964 95200
rect 151904 94694 152106 94754
rect 151678 94150 151828 94210
rect 151678 92445 151738 94150
rect 152046 92445 152106 94694
rect 151675 92444 151741 92445
rect 151675 92380 151676 92444
rect 151740 92380 151741 92444
rect 151675 92379 151741 92380
rect 152043 92444 152109 92445
rect 152043 92380 152044 92444
rect 152108 92380 152109 92444
rect 152043 92379 152109 92380
rect 151123 91492 151189 91493
rect 151123 91428 151124 91492
rect 151188 91428 151189 91492
rect 151123 91427 151189 91428
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 82894 153854 93100
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 86614 157574 93100
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 93100
rect 166214 88229 166274 135491
rect 166950 115837 167010 271899
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 167514 169174 168134 204618
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 167514 133174 168134 168618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 168971 142220 169037 142221
rect 168971 142156 168972 142220
rect 169036 142156 169037 142220
rect 168971 142155 169037 142156
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 166947 115836 167013 115837
rect 166947 115772 166948 115836
rect 167012 115772 167013 115836
rect 166947 115771 167013 115772
rect 166947 98020 167013 98021
rect 166947 97956 166948 98020
rect 167012 97956 167013 98020
rect 166947 97955 167013 97956
rect 166395 97204 166461 97205
rect 166395 97140 166396 97204
rect 166460 97140 166461 97204
rect 166395 97139 166461 97140
rect 166398 92309 166458 97139
rect 166950 95165 167010 97955
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 166947 95164 167013 95165
rect 166947 95100 166948 95164
rect 167012 95100 167013 95164
rect 166947 95099 167013 95100
rect 166395 92308 166461 92309
rect 166395 92244 166396 92308
rect 166460 92244 166461 92308
rect 166395 92243 166461 92244
rect 166211 88228 166277 88229
rect 166211 88164 166212 88228
rect 166276 88164 166277 88228
rect 166211 88163 166277 88164
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 61174 168134 96618
rect 168974 89725 169034 142155
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 170259 128620 170325 128621
rect 170259 128556 170260 128620
rect 170324 128556 170325 128620
rect 170259 128555 170325 128556
rect 169155 127124 169221 127125
rect 169155 127060 169156 127124
rect 169220 127060 169221 127124
rect 169155 127059 169221 127060
rect 168971 89724 169037 89725
rect 168971 89660 168972 89724
rect 169036 89660 169037 89724
rect 168971 89659 169037 89660
rect 169158 78573 169218 127059
rect 170262 80069 170322 128555
rect 170443 102236 170509 102237
rect 170443 102172 170444 102236
rect 170508 102172 170509 102236
rect 170443 102171 170509 102172
rect 170446 91085 170506 102171
rect 171234 100894 171854 136338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 173019 127260 173085 127261
rect 173019 127196 173020 127260
rect 173084 127196 173085 127260
rect 173019 127195 173085 127196
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 170443 91084 170509 91085
rect 170443 91020 170444 91084
rect 170508 91020 170509 91084
rect 170443 91019 170509 91020
rect 170259 80068 170325 80069
rect 170259 80004 170260 80068
rect 170324 80004 170325 80068
rect 170259 80003 170325 80004
rect 169155 78572 169221 78573
rect 169155 78508 169156 78572
rect 169220 78508 169221 78572
rect 169155 78507 169221 78508
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 64894 171854 100338
rect 173022 81429 173082 127195
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 173019 81428 173085 81429
rect 173019 81364 173020 81428
rect 173084 81364 173085 81428
rect 173019 81363 173085 81364
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 277174 204134 312618
rect 203514 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 204134 277174
rect 203514 276854 204134 276938
rect 203514 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 204134 276854
rect 203514 241174 204134 276618
rect 203514 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 204134 241174
rect 203514 240854 204134 240938
rect 203514 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 204134 240854
rect 203514 205174 204134 240618
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 280894 207854 316338
rect 207234 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 207854 280894
rect 207234 280574 207854 280658
rect 207234 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 207854 280574
rect 207234 244894 207854 280338
rect 207234 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 207854 244894
rect 207234 244574 207854 244658
rect 207234 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 207854 244574
rect 207234 208894 207854 244338
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 284614 211574 320058
rect 210954 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 211574 284614
rect 210954 284294 211574 284378
rect 210954 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 211574 284294
rect 210954 248614 211574 284058
rect 210954 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 211574 248614
rect 210954 248294 211574 248378
rect 210954 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 211574 248294
rect 210954 212614 211574 248058
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 178000 218414 182898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 223174 222134 258618
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 178000 222134 186618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 262894 225854 298338
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 226894 225854 262338
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 178000 225854 190338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 266614 229574 302058
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228954 230614 229574 266058
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 178000 229574 194058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 178000 236414 200898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385174 240134 420618
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 349174 240134 384618
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 239514 313174 240134 348618
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 239514 277174 240134 312618
rect 239514 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 240134 277174
rect 239514 276854 240134 276938
rect 239514 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 240134 276854
rect 239514 241174 240134 276618
rect 239514 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 240134 241174
rect 239514 240854 240134 240938
rect 239514 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 240134 240854
rect 239514 205174 240134 240618
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 239514 178000 240134 204618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 352894 243854 388338
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 243234 316894 243854 352338
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 243234 280894 243854 316338
rect 243234 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 243854 280894
rect 243234 280574 243854 280658
rect 243234 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 243854 280574
rect 243234 244894 243854 280338
rect 243234 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 243854 244894
rect 243234 244574 243854 244658
rect 243234 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 243854 244574
rect 243234 208894 243854 244338
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 243234 178000 243854 208338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 356614 247574 392058
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 246954 320614 247574 356058
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 246954 284614 247574 320058
rect 246954 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 247574 284614
rect 246954 284294 247574 284378
rect 246954 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 247574 284294
rect 246954 248614 247574 284058
rect 246954 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 247574 248614
rect 246954 248294 247574 248378
rect 246954 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 247574 248294
rect 246954 212614 247574 248058
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 246954 178000 247574 212058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 254531 296852 254597 296853
rect 254531 296788 254532 296852
rect 254596 296788 254597 296852
rect 254531 296787 254597 296788
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 249379 177308 249445 177309
rect 249379 177244 249380 177308
rect 249444 177244 249445 177308
rect 249379 177243 249445 177244
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 140614 211574 176058
rect 249195 176084 249261 176085
rect 249195 176020 249196 176084
rect 249260 176020 249261 176084
rect 249195 176019 249261 176020
rect 249198 174317 249258 176019
rect 249195 174316 249261 174317
rect 249195 174252 249196 174316
rect 249260 174252 249261 174316
rect 249195 174251 249261 174252
rect 249382 173365 249442 177243
rect 249379 173364 249445 173365
rect 249379 173300 249380 173364
rect 249444 173300 249445 173364
rect 249379 173299 249445 173300
rect 227874 165454 228194 165486
rect 227874 165218 227916 165454
rect 228152 165218 228194 165454
rect 227874 165134 228194 165218
rect 227874 164898 227916 165134
rect 228152 164898 228194 165134
rect 227874 164866 228194 164898
rect 237805 165454 238125 165486
rect 237805 165218 237847 165454
rect 238083 165218 238125 165454
rect 237805 165134 238125 165218
rect 237805 164898 237847 165134
rect 238083 164898 238125 165134
rect 237805 164866 238125 164898
rect 251771 148204 251837 148205
rect 251771 148140 251772 148204
rect 251836 148140 251837 148204
rect 251771 148139 251837 148140
rect 222910 147454 223230 147486
rect 222910 147218 222952 147454
rect 223188 147218 223230 147454
rect 222910 147134 223230 147218
rect 222910 146898 222952 147134
rect 223188 146898 223230 147134
rect 222910 146866 223230 146898
rect 232840 147454 233160 147486
rect 232840 147218 232882 147454
rect 233118 147218 233160 147454
rect 232840 147134 233160 147218
rect 232840 146898 232882 147134
rect 233118 146898 233160 147134
rect 232840 146866 233160 146898
rect 242771 147454 243091 147486
rect 242771 147218 242813 147454
rect 243049 147218 243091 147454
rect 242771 147134 243091 147218
rect 242771 146898 242813 147134
rect 243049 146898 243091 147134
rect 242771 146866 243091 146898
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 227874 129454 228194 129486
rect 227874 129218 227916 129454
rect 228152 129218 228194 129454
rect 227874 129134 228194 129218
rect 227874 128898 227916 129134
rect 228152 128898 228194 129134
rect 227874 128866 228194 128898
rect 237805 129454 238125 129486
rect 237805 129218 237847 129454
rect 238083 129218 238125 129454
rect 237805 129134 238125 129218
rect 237805 128898 237847 129134
rect 238083 128898 238125 129134
rect 237805 128866 238125 128898
rect 251774 112709 251834 148139
rect 253794 147454 254414 182898
rect 254534 163437 254594 296787
rect 257514 295174 258134 330618
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 223174 258134 258618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 261234 298894 261854 334338
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 261234 262894 261854 298338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264954 302614 265574 338058
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 263547 269244 263613 269245
rect 263547 269180 263548 269244
rect 263612 269180 263613 269244
rect 263547 269179 263613 269180
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 258395 245716 258461 245717
rect 258395 245652 258396 245716
rect 258460 245652 258461 245716
rect 258395 245651 258461 245652
rect 258398 238770 258458 245651
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 256739 185604 256805 185605
rect 256739 185540 256740 185604
rect 256804 185540 256805 185604
rect 256739 185539 256805 185540
rect 255267 178804 255333 178805
rect 255267 178740 255268 178804
rect 255332 178740 255333 178804
rect 255267 178739 255333 178740
rect 254531 163436 254597 163437
rect 254531 163372 254532 163436
rect 254596 163372 254597 163436
rect 254531 163371 254597 163372
rect 255270 147525 255330 178739
rect 255267 147524 255333 147525
rect 255267 147460 255268 147524
rect 255332 147460 255333 147524
rect 255267 147459 255333 147460
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 251955 142356 252021 142357
rect 251955 142292 251956 142356
rect 252020 142292 252021 142356
rect 251955 142291 252021 142292
rect 251958 130933 252018 142291
rect 251955 130932 252021 130933
rect 251955 130868 251956 130932
rect 252020 130868 252021 130932
rect 251955 130867 252021 130868
rect 251771 112708 251837 112709
rect 251771 112644 251772 112708
rect 251836 112644 251837 112708
rect 251771 112643 251837 112644
rect 222910 111454 223230 111486
rect 222910 111218 222952 111454
rect 223188 111218 223230 111454
rect 222910 111134 223230 111218
rect 222910 110898 222952 111134
rect 223188 110898 223230 111134
rect 222910 110866 223230 110898
rect 232840 111454 233160 111486
rect 232840 111218 232882 111454
rect 233118 111218 233160 111454
rect 232840 111134 233160 111218
rect 232840 110898 232882 111134
rect 233118 110898 233160 111134
rect 232840 110866 233160 110898
rect 242771 111454 243091 111486
rect 242771 111218 242813 111454
rect 243049 111218 243091 111454
rect 242771 111134 243091 111218
rect 242771 110898 242813 111134
rect 243049 110898 243091 111134
rect 242771 110866 243091 110898
rect 253794 111454 254414 146898
rect 256742 140453 256802 185539
rect 257514 151174 258134 186618
rect 258214 238710 258458 238770
rect 258214 151830 258274 238710
rect 261234 226894 261854 262338
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 190894 261854 226338
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 258395 177580 258461 177581
rect 258395 177516 258396 177580
rect 258460 177516 258461 177580
rect 258395 177515 258461 177516
rect 258398 155277 258458 177515
rect 259499 177444 259565 177445
rect 259499 177380 259500 177444
rect 259564 177380 259565 177444
rect 259499 177379 259565 177380
rect 259502 160853 259562 177379
rect 260051 176764 260117 176765
rect 260051 176700 260052 176764
rect 260116 176700 260117 176764
rect 260051 176699 260117 176700
rect 259499 160852 259565 160853
rect 259499 160788 259500 160852
rect 259564 160788 259565 160852
rect 259499 160787 259565 160788
rect 258395 155276 258461 155277
rect 258395 155212 258396 155276
rect 258460 155212 258461 155276
rect 258395 155211 258461 155212
rect 258579 153508 258645 153509
rect 258579 153444 258580 153508
rect 258644 153444 258645 153508
rect 258579 153443 258645 153444
rect 258214 151770 258458 151830
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 256739 140452 256805 140453
rect 256739 140388 256740 140452
rect 256804 140388 256805 140452
rect 256739 140387 256805 140388
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 214419 105228 214485 105229
rect 214419 105164 214420 105228
rect 214484 105164 214485 105228
rect 214419 105163 214485 105164
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 214422 93805 214482 105163
rect 214419 93804 214485 93805
rect 214419 93740 214420 93804
rect 214484 93740 214485 93804
rect 214419 93739 214485 93740
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 75454 218414 94000
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 79174 222134 94000
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 82894 225854 94000
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 86614 229574 94000
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 93454 236414 94000
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 61174 240134 94000
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 64894 243854 94000
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 68614 247574 94000
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 115174 258134 150618
rect 258398 146301 258458 151770
rect 258395 146300 258461 146301
rect 258395 146236 258396 146300
rect 258460 146236 258461 146300
rect 258395 146235 258461 146236
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 258582 112981 258642 153443
rect 258579 112980 258645 112981
rect 258579 112916 258580 112980
rect 258644 112916 258645 112980
rect 258579 112915 258645 112916
rect 260054 96661 260114 176699
rect 260971 175948 261037 175949
rect 260971 175884 260972 175948
rect 261036 175884 261037 175948
rect 260971 175883 261037 175884
rect 260974 170373 261034 175883
rect 260971 170372 261037 170373
rect 260971 170308 260972 170372
rect 261036 170308 261037 170372
rect 260971 170307 261037 170308
rect 261234 154894 261854 190338
rect 262811 175404 262877 175405
rect 262811 175340 262812 175404
rect 262876 175340 262877 175404
rect 262811 175339 262877 175340
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 260051 96660 260117 96661
rect 260051 96596 260052 96660
rect 260116 96596 260117 96660
rect 260051 96595 260117 96596
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 82894 261854 118338
rect 262814 96797 262874 175339
rect 263550 144533 263610 269179
rect 264954 266614 265574 302058
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 230614 265574 266058
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 267779 218652 267845 218653
rect 267779 218588 267780 218652
rect 267844 218588 267845 218652
rect 267779 218587 267845 218588
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 263731 191044 263797 191045
rect 263731 190980 263732 191044
rect 263796 190980 263797 191044
rect 263731 190979 263797 190980
rect 263547 144532 263613 144533
rect 263547 144468 263548 144532
rect 263612 144468 263613 144532
rect 263547 144467 263613 144468
rect 263734 138821 263794 190979
rect 264954 158614 265574 194058
rect 266307 192540 266373 192541
rect 266307 192476 266308 192540
rect 266372 192476 266373 192540
rect 266307 192475 266373 192476
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 263731 138820 263797 138821
rect 263731 138756 263732 138820
rect 263796 138756 263797 138820
rect 263731 138755 263797 138756
rect 264954 122614 265574 158058
rect 266310 153373 266370 192475
rect 266307 153372 266373 153373
rect 266307 153308 266308 153372
rect 266372 153308 266373 153372
rect 266307 153307 266373 153308
rect 267782 140861 267842 218587
rect 269067 203556 269133 203557
rect 269067 203492 269068 203556
rect 269132 203492 269133 203556
rect 269067 203491 269133 203492
rect 269070 157453 269130 203491
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 269067 157452 269133 157453
rect 269067 157388 269068 157452
rect 269132 157388 269133 157452
rect 269067 157387 269133 157388
rect 267779 140860 267845 140861
rect 267779 140796 267780 140860
rect 267844 140796 267845 140860
rect 267779 140795 267845 140796
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 262811 96796 262877 96797
rect 262811 96732 262812 96796
rect 262876 96732 262877 96796
rect 262811 96731 262877 96732
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 349174 276134 384618
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 277174 276134 312618
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 205174 276134 240618
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 169174 276134 204618
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 133174 276134 168618
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 352894 279854 388338
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 280894 279854 316338
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279234 172894 279854 208338
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 279234 136894 279854 172338
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 100894 279854 136338
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 356614 283574 392058
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 282954 284614 283574 320058
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 282954 248614 283574 284058
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 282954 176614 283574 212058
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 178000 308414 200898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 178000 312134 204618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 178000 315854 208338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 320219 225588 320285 225589
rect 320219 225524 320220 225588
rect 320284 225524 320285 225588
rect 320219 225523 320285 225524
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 178000 319574 212058
rect 320222 190470 320282 225523
rect 325794 219454 326414 254898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 331259 300932 331325 300933
rect 331259 300868 331260 300932
rect 331324 300868 331325 300932
rect 331259 300867 331325 300868
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 327027 222868 327093 222869
rect 327027 222804 327028 222868
rect 327092 222804 327093 222868
rect 327027 222803 327093 222804
rect 329514 222854 330134 222938
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 324267 196620 324333 196621
rect 324267 196556 324268 196620
rect 324332 196556 324333 196620
rect 324267 196555 324333 196556
rect 320222 190410 321386 190470
rect 321326 170645 321386 190410
rect 321323 170644 321389 170645
rect 321323 170580 321324 170644
rect 321388 170580 321389 170644
rect 321323 170579 321389 170580
rect 314208 165454 314528 165486
rect 314208 165218 314250 165454
rect 314486 165218 314528 165454
rect 314208 165134 314528 165218
rect 314208 164898 314250 165134
rect 314486 164898 314528 165134
rect 314208 164866 314528 164898
rect 317472 165454 317792 165486
rect 317472 165218 317514 165454
rect 317750 165218 317792 165454
rect 317472 165134 317792 165218
rect 317472 164898 317514 165134
rect 317750 164898 317792 165134
rect 317472 164866 317792 164898
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 312576 147454 312896 147486
rect 312576 147218 312618 147454
rect 312854 147218 312896 147454
rect 312576 147134 312896 147218
rect 312576 146898 312618 147134
rect 312854 146898 312896 147134
rect 312576 146866 312896 146898
rect 315840 147454 316160 147486
rect 315840 147218 315882 147454
rect 316118 147218 316160 147454
rect 315840 147134 316160 147218
rect 315840 146898 315882 147134
rect 316118 146898 316160 147134
rect 315840 146866 316160 146898
rect 319104 147454 319424 147486
rect 319104 147218 319146 147454
rect 319382 147218 319424 147454
rect 319104 147134 319424 147218
rect 319104 146898 319146 147134
rect 319382 146898 319424 147134
rect 319104 146866 319424 146898
rect 307707 146436 307773 146437
rect 307707 146372 307708 146436
rect 307772 146372 307773 146436
rect 307707 146371 307773 146372
rect 307710 145621 307770 146371
rect 307707 145620 307773 145621
rect 307707 145556 307708 145620
rect 307772 145556 307773 145620
rect 307707 145555 307773 145556
rect 302739 134060 302805 134061
rect 302739 133996 302740 134060
rect 302804 133996 302805 134060
rect 302739 133995 302805 133996
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 299979 118148 300045 118149
rect 299979 118084 299980 118148
rect 300044 118084 300045 118148
rect 299979 118083 300045 118084
rect 298691 97748 298757 97749
rect 298691 97684 298692 97748
rect 298756 97684 298757 97748
rect 298691 97683 298757 97684
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 298694 57221 298754 97683
rect 298691 57220 298757 57221
rect 298691 57156 298692 57220
rect 298756 57156 298757 57220
rect 298691 57155 298757 57156
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 299982 30973 300042 118083
rect 300954 86614 301574 122058
rect 301819 113524 301885 113525
rect 301819 113460 301820 113524
rect 301884 113460 301885 113524
rect 301819 113459 301885 113460
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 301822 54501 301882 113459
rect 301819 54500 301885 54501
rect 301819 54436 301820 54500
rect 301884 54436 301885 54500
rect 301819 54435 301885 54436
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 299979 30972 300045 30973
rect 299979 30908 299980 30972
rect 300044 30908 300045 30972
rect 299979 30907 300045 30908
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 14614 301574 50058
rect 302742 29613 302802 133995
rect 305499 130116 305565 130117
rect 305499 130052 305500 130116
rect 305564 130052 305565 130116
rect 305499 130051 305565 130052
rect 302923 112164 302989 112165
rect 302923 112100 302924 112164
rect 302988 112100 302989 112164
rect 302923 112099 302989 112100
rect 302926 61437 302986 112099
rect 304211 104140 304277 104141
rect 304211 104076 304212 104140
rect 304276 104076 304277 104140
rect 304211 104075 304277 104076
rect 302923 61436 302989 61437
rect 302923 61372 302924 61436
rect 302988 61372 302989 61436
rect 302923 61371 302989 61372
rect 302739 29612 302805 29613
rect 302739 29548 302740 29612
rect 302804 29548 302805 29612
rect 302739 29547 302805 29548
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 304214 13021 304274 104075
rect 304395 101964 304461 101965
rect 304395 101900 304396 101964
rect 304460 101900 304461 101964
rect 304395 101899 304461 101900
rect 304398 62797 304458 101899
rect 304395 62796 304461 62797
rect 304395 62732 304396 62796
rect 304460 62732 304461 62796
rect 304395 62731 304461 62732
rect 305502 47565 305562 130051
rect 314208 129454 314528 129486
rect 314208 129218 314250 129454
rect 314486 129218 314528 129454
rect 314208 129134 314528 129218
rect 314208 128898 314250 129134
rect 314486 128898 314528 129134
rect 314208 128866 314528 128898
rect 317472 129454 317792 129486
rect 317472 129218 317514 129454
rect 317750 129218 317792 129454
rect 317472 129134 317792 129218
rect 317472 128898 317514 129134
rect 317750 128898 317792 129134
rect 317472 128866 317792 128898
rect 307155 114068 307221 114069
rect 307155 114004 307156 114068
rect 307220 114004 307221 114068
rect 307155 114003 307221 114004
rect 305683 99652 305749 99653
rect 305683 99588 305684 99652
rect 305748 99588 305749 99652
rect 305683 99587 305749 99588
rect 305499 47564 305565 47565
rect 305499 47500 305500 47564
rect 305564 47500 305565 47564
rect 305499 47499 305565 47500
rect 305686 18597 305746 99587
rect 306971 97068 307037 97069
rect 306971 97004 306972 97068
rect 307036 97004 307037 97068
rect 306971 97003 307037 97004
rect 305683 18596 305749 18597
rect 305683 18532 305684 18596
rect 305748 18532 305749 18596
rect 305683 18531 305749 18532
rect 304211 13020 304277 13021
rect 304211 12956 304212 13020
rect 304276 12956 304277 13020
rect 304211 12955 304277 12956
rect 306974 4861 307034 97003
rect 307158 32469 307218 114003
rect 312576 111454 312896 111486
rect 312576 111218 312618 111454
rect 312854 111218 312896 111454
rect 312576 111134 312896 111218
rect 312576 110898 312618 111134
rect 312854 110898 312896 111134
rect 312576 110866 312896 110898
rect 315840 111454 316160 111486
rect 315840 111218 315882 111454
rect 316118 111218 316160 111454
rect 315840 111134 316160 111218
rect 315840 110898 315882 111134
rect 316118 110898 316160 111134
rect 315840 110866 316160 110898
rect 319104 111454 319424 111486
rect 319104 111218 319146 111454
rect 319382 111218 319424 111454
rect 319104 111134 319424 111218
rect 319104 110898 319146 111134
rect 319382 110898 319424 111134
rect 319104 110866 319424 110898
rect 324270 100877 324330 196555
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 324267 100876 324333 100877
rect 324267 100812 324268 100876
rect 324332 100812 324333 100876
rect 324267 100811 324333 100812
rect 307794 93454 308414 94000
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307155 32468 307221 32469
rect 307155 32404 307156 32468
rect 307220 32404 307221 32468
rect 307155 32403 307221 32404
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 306971 4860 307037 4861
rect 306971 4796 306972 4860
rect 307036 4796 307037 4860
rect 306971 4795 307037 4796
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 61174 312134 94000
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 64894 315854 94000
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 68614 319574 94000
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 75454 326414 110898
rect 327030 106317 327090 222803
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 327211 213212 327277 213213
rect 327211 213148 327212 213212
rect 327276 213148 327277 213212
rect 327211 213147 327277 213148
rect 327214 107813 327274 213147
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 327211 107812 327277 107813
rect 327211 107748 327212 107812
rect 327276 107748 327277 107812
rect 327211 107747 327277 107748
rect 327027 106316 327093 106317
rect 327027 106252 327028 106316
rect 327092 106252 327093 106316
rect 327027 106251 327093 106252
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 79174 330134 114618
rect 331262 98157 331322 300867
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 335123 291956 335189 291957
rect 335123 291892 335124 291956
rect 335188 291892 335189 291956
rect 335123 291891 335189 291892
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 334019 210356 334085 210357
rect 334019 210292 334020 210356
rect 334084 210292 334085 210356
rect 334019 210291 334085 210292
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 332547 178804 332613 178805
rect 332547 178740 332548 178804
rect 332612 178740 332613 178804
rect 332547 178739 332613 178740
rect 331443 177308 331509 177309
rect 331443 177244 331444 177308
rect 331508 177244 331509 177308
rect 331443 177243 331509 177244
rect 331446 114749 331506 177243
rect 331443 114748 331509 114749
rect 331443 114684 331444 114748
rect 331508 114684 331509 114748
rect 331443 114683 331509 114684
rect 332550 110669 332610 178739
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 332547 110668 332613 110669
rect 332547 110604 332548 110668
rect 332612 110604 332613 110668
rect 332547 110603 332613 110604
rect 331259 98156 331325 98157
rect 331259 98092 331260 98156
rect 331324 98092 331325 98156
rect 331259 98091 331325 98092
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 82894 333854 118338
rect 334022 101013 334082 210291
rect 334203 178940 334269 178941
rect 334203 178876 334204 178940
rect 334268 178876 334269 178940
rect 334203 178875 334269 178876
rect 334206 109581 334266 178875
rect 334203 109580 334269 109581
rect 334203 109516 334204 109580
rect 334268 109516 334269 109580
rect 334203 109515 334269 109516
rect 335126 109173 335186 291891
rect 336954 266614 337574 302058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 342115 291276 342181 291277
rect 342115 291212 342116 291276
rect 342180 291212 342181 291276
rect 342115 291211 342181 291212
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 340091 264212 340157 264213
rect 340091 264148 340092 264212
rect 340156 264148 340157 264212
rect 340091 264147 340157 264148
rect 338619 259588 338685 259589
rect 338619 259524 338620 259588
rect 338684 259524 338685 259588
rect 338619 259523 338685 259524
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336779 194580 336845 194581
rect 336779 194516 336780 194580
rect 336844 194516 336845 194580
rect 336779 194515 336845 194516
rect 335491 180028 335557 180029
rect 335491 179964 335492 180028
rect 335556 179964 335557 180028
rect 335491 179963 335557 179964
rect 335494 115973 335554 179963
rect 336782 135285 336842 194515
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 338251 179348 338317 179349
rect 338251 179284 338252 179348
rect 338316 179284 338317 179348
rect 338251 179283 338317 179284
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336779 135284 336845 135285
rect 336779 135220 336780 135284
rect 336844 135220 336845 135284
rect 336779 135219 336845 135220
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 335491 115972 335557 115973
rect 335491 115908 335492 115972
rect 335556 115908 335557 115972
rect 335491 115907 335557 115908
rect 335123 109172 335189 109173
rect 335123 109108 335124 109172
rect 335188 109108 335189 109172
rect 335123 109107 335189 109108
rect 334019 101012 334085 101013
rect 334019 100948 334020 101012
rect 334084 100948 334085 101012
rect 334019 100947 334085 100948
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 86614 337574 122058
rect 338254 110533 338314 179283
rect 338622 165749 338682 259523
rect 338619 165748 338685 165749
rect 338619 165684 338620 165748
rect 338684 165684 338685 165748
rect 338619 165683 338685 165684
rect 338251 110532 338317 110533
rect 338251 110468 338252 110532
rect 338316 110468 338317 110532
rect 338251 110467 338317 110468
rect 340094 99517 340154 264147
rect 342118 138141 342178 291211
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 342299 211852 342365 211853
rect 342299 211788 342300 211852
rect 342364 211788 342365 211852
rect 342299 211787 342365 211788
rect 342115 138140 342181 138141
rect 342115 138076 342116 138140
rect 342180 138076 342181 138140
rect 342115 138075 342181 138076
rect 342302 106453 342362 211787
rect 343794 201454 344414 236898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 345059 236604 345125 236605
rect 345059 236540 345060 236604
rect 345124 236540 345125 236604
rect 345059 236539 345125 236540
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 342299 106452 342365 106453
rect 342299 106388 342300 106452
rect 342364 106388 342365 106452
rect 342299 106387 342365 106388
rect 340091 99516 340157 99517
rect 340091 99452 340092 99516
rect 340156 99452 340157 99516
rect 340091 99451 340157 99452
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 93454 344414 128898
rect 345062 114613 345122 236539
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 345059 114612 345125 114613
rect 345059 114548 345060 114612
rect 345124 114548 345125 114612
rect 345059 114547 345125 114548
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 89610 273218 89846 273454
rect 89610 272898 89846 273134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 74250 255218 74486 255454
rect 74250 254898 74486 255134
rect 104970 255218 105206 255454
rect 104970 254898 105206 255134
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 69128 165218 69364 165454
rect 69128 164898 69364 165134
rect 164192 165218 164428 165454
rect 164192 164898 164428 165134
rect 69808 147218 70044 147454
rect 69808 146898 70044 147134
rect 163512 147218 163748 147454
rect 163512 146898 163748 147134
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 69128 129218 69364 129454
rect 69128 128898 69364 129134
rect 164192 129218 164428 129454
rect 164192 128898 164428 129134
rect 69808 111218 70044 111454
rect 69808 110898 70044 111134
rect 163512 111218 163748 111454
rect 163512 110898 163748 111134
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 203546 276938 203782 277174
rect 203866 276938 204102 277174
rect 203546 276618 203782 276854
rect 203866 276618 204102 276854
rect 203546 240938 203782 241174
rect 203866 240938 204102 241174
rect 203546 240618 203782 240854
rect 203866 240618 204102 240854
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 207266 280658 207502 280894
rect 207586 280658 207822 280894
rect 207266 280338 207502 280574
rect 207586 280338 207822 280574
rect 207266 244658 207502 244894
rect 207586 244658 207822 244894
rect 207266 244338 207502 244574
rect 207586 244338 207822 244574
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 210986 284378 211222 284614
rect 211306 284378 211542 284614
rect 210986 284058 211222 284294
rect 211306 284058 211542 284294
rect 210986 248378 211222 248614
rect 211306 248378 211542 248614
rect 210986 248058 211222 248294
rect 211306 248058 211542 248294
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 239546 276938 239782 277174
rect 239866 276938 240102 277174
rect 239546 276618 239782 276854
rect 239866 276618 240102 276854
rect 239546 240938 239782 241174
rect 239866 240938 240102 241174
rect 239546 240618 239782 240854
rect 239866 240618 240102 240854
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 243266 280658 243502 280894
rect 243586 280658 243822 280894
rect 243266 280338 243502 280574
rect 243586 280338 243822 280574
rect 243266 244658 243502 244894
rect 243586 244658 243822 244894
rect 243266 244338 243502 244574
rect 243586 244338 243822 244574
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 246986 284378 247222 284614
rect 247306 284378 247542 284614
rect 246986 284058 247222 284294
rect 247306 284058 247542 284294
rect 246986 248378 247222 248614
rect 247306 248378 247542 248614
rect 246986 248058 247222 248294
rect 247306 248058 247542 248294
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 227916 165218 228152 165454
rect 227916 164898 228152 165134
rect 237847 165218 238083 165454
rect 237847 164898 238083 165134
rect 222952 147218 223188 147454
rect 222952 146898 223188 147134
rect 232882 147218 233118 147454
rect 232882 146898 233118 147134
rect 242813 147218 243049 147454
rect 242813 146898 243049 147134
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 227916 129218 228152 129454
rect 227916 128898 228152 129134
rect 237847 129218 238083 129454
rect 237847 128898 238083 129134
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 222952 111218 223188 111454
rect 222952 110898 223188 111134
rect 232882 111218 233118 111454
rect 232882 110898 233118 111134
rect 242813 111218 243049 111454
rect 242813 110898 243049 111134
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 314250 165218 314486 165454
rect 314250 164898 314486 165134
rect 317514 165218 317750 165454
rect 317514 164898 317750 165134
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 312618 147218 312854 147454
rect 312618 146898 312854 147134
rect 315882 147218 316118 147454
rect 315882 146898 316118 147134
rect 319146 147218 319382 147454
rect 319146 146898 319382 147134
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 314250 129218 314486 129454
rect 314250 128898 314486 129134
rect 317514 129218 317750 129454
rect 317514 128898 317750 129134
rect 312618 111218 312854 111454
rect 312618 110898 312854 111134
rect 315882 111218 316118 111454
rect 315882 110898 316118 111134
rect 319146 111218 319382 111454
rect 319146 110898 319382 111134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 89610 273454
rect 89846 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 89610 273134
rect 89846 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 74250 255454
rect 74486 255218 104970 255454
rect 105206 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 74250 255134
rect 74486 254898 104970 255134
rect 105206 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 69128 165454
rect 69364 165218 164192 165454
rect 164428 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 227916 165454
rect 228152 165218 237847 165454
rect 238083 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 314250 165454
rect 314486 165218 317514 165454
rect 317750 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 69128 165134
rect 69364 164898 164192 165134
rect 164428 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 227916 165134
rect 228152 164898 237847 165134
rect 238083 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 314250 165134
rect 314486 164898 317514 165134
rect 317750 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 69808 147454
rect 70044 147218 163512 147454
rect 163748 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 222952 147454
rect 223188 147218 232882 147454
rect 233118 147218 242813 147454
rect 243049 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 312618 147454
rect 312854 147218 315882 147454
rect 316118 147218 319146 147454
rect 319382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 69808 147134
rect 70044 146898 163512 147134
rect 163748 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 222952 147134
rect 223188 146898 232882 147134
rect 233118 146898 242813 147134
rect 243049 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 312618 147134
rect 312854 146898 315882 147134
rect 316118 146898 319146 147134
rect 319382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 69128 129454
rect 69364 129218 164192 129454
rect 164428 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 227916 129454
rect 228152 129218 237847 129454
rect 238083 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 314250 129454
rect 314486 129218 317514 129454
rect 317750 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 69128 129134
rect 69364 128898 164192 129134
rect 164428 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 227916 129134
rect 228152 128898 237847 129134
rect 238083 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 314250 129134
rect 314486 128898 317514 129134
rect 317750 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 69808 111454
rect 70044 111218 163512 111454
rect 163748 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 222952 111454
rect 223188 111218 232882 111454
rect 233118 111218 242813 111454
rect 243049 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 312618 111454
rect 312854 111218 315882 111454
rect 316118 111218 319146 111454
rect 319382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 69808 111134
rect 70044 110898 163512 111134
rect 163748 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 222952 111134
rect 223188 110898 232882 111134
rect 233118 110898 242813 111134
rect 243049 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 312618 111134
rect 312854 110898 315882 111134
rect 316118 110898 319146 111134
rect 319382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_1kbyte_1rw1r_32x256_8  openram_1kB
timestamp 0
transform 1 0 68800 0 1 95100
box 0 0 95956 79500
use wb_bridge_2way  wb_bridge_2way
timestamp 0
transform 1 0 310000 0 1 96000
box 0 144 12000 80000
use wb_openram_wrapper  wb_openram_wrapper
timestamp 0
transform 1 0 217000 0 1 96000
box 0 144 32000 79688
use wrapped_function_generator  wrapped_function_generator_0
timestamp 0
transform 1 0 70000 0 1 240000
box 0 0 50000 52000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 94000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 176600 74414 238000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 176600 110414 238000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 294000 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 294000 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 176600 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 178000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 94000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 176600 78134 238000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 176600 114134 238000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 294000 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 294000 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 176600 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 178000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 94000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 176600 81854 238000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 176600 117854 238000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 294000 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 294000 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 176600 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 178000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 94000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 176600 85574 238000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 176600 121574 238000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 294000 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 294000 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 176600 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 178000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 94000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 94000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 176600 99854 238000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 294000 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 176600 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 178000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 178000 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 94000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 94000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 176600 103574 238000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 176600 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 294000 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 176600 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 178000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 178000 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 94000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 94000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 176600 92414 238000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 294000 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 176600 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 176600 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 178000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 178000 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 94000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 94000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 176600 96134 238000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 294000 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 176600 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 178000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 178000 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
